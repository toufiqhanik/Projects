.Option brief ingold=2 accurate
.OPTION MEASDGT=8
.OPTION NUMDGT=10
+ RUNLVL=5 ACCURATE
.op

.PARAM VDD_VALUE= 1.2
.PARAM VDD_HALF= 0.6
.OPTION BRIEF=1

.OPTION POST=2
.OPTION MEASFORM=3
.OPTION PROBE=1

******
.PARAM vth_pmos_pv=GAUSS(-0.3021,0.1,1)
.PARAM vth_nmos_pv=GAUSS(0.322,0.1,1)
.PARAM toxm_pmos_pv=GAUSS(1.26E-009,0.01,1)
.PARAM toxm_nmos_pv=GAUSS(1.14E-09,0.01,1)
.PARAM LMIN_pv=GAUSS(50E-09,0.1,3)

******

VSUPPLY VDD 0 VDD_VALUE
VSUPPLYGND GND 0 0

Vinputclk CLK GND PWL (0 0 136.9n 0 137n VDD_VALUE 150n VDD_VALUE)

Vinputrst reset GND PWL(0 VDD_VALUE 1.9n VDD_VALUE 2n 0 2.9n 0 3n VDD_VALUE)
*depending on the delay of buffer ro_control should be changed


.TRAN 138N 150N START=0N SWEEP MONTE=5 FIRSTRUN =1

.include './trans_model_nk'
.temp tempvar

******** NAND MODEL ***********
* The subcircuit for NAND
.SUBCKT NAND2_X1
+ A1 A2
+ ZN
+ VDDx GNDx
M_i_1 net_0 A1 GNDx GNDx NMOS_VTL_pv W=0.415000U L='LMIN_pv'
M_i_0 ZN A2 net_0 GNDx NMOS_VTL_pv W=0.415000U L='LMIN_pv'
M_i_11 ZN A2 VDDx VDDx PMOS_VTL_pv W=0.630000U L='LMIN_pv'
M_i_10 VDDx A1 ZN VDDx PMOS_VTL_pv W=0.630000U L='LMIN_pv'
.ENDS

******** INV MODEL ***********
* The subcircuit for INV
.SUBCKT INV_X1
+ A1
+ ZN
+ VDDx GNDx
M_i_0 ZN A1 GNDx GNDx NMOS_VTL_pv W=0.415000U L='LMIN_pv'
M_i_10 ZN A1 VDDx VDDx PMOS_VTL_pv W=0.630000U L='LMIN_pv'
.ENDS

******** DFFR_X1 MODEL ***********
* The subcircuit for DFFR_X1
.SUBCKT DFFR_X1
+ D CK RN
+ Q QN
+ VDDx GNDx

*.PININFO D:I RN:I CK:I Q:O QN:O VDDx:P GNDx:G 
M_i_0 GNDx CK net_000 GNDx NMOS_VTL_pv W=0.210000U L='LMIN_pv'
M_i_7 net_001 net_000 GNDx GNDx NMOS_VTL_pv W=0.210000U L='LMIN_pv'
M_i_13 net_002 D GNDx GNDx NMOS_VTL_pv W=0.275000U L='LMIN_pv'
M_i_18 net_003 net_000 net_002 GNDx NMOS_VTL_pv W=0.275000U L='LMIN_pv'
M_i_24 net_004 net_001 net_003 GNDx NMOS_VTL_pv W=0.090000U L='LMIN_pv'
M_i_28 net_005 net_006 net_004 GNDx NMOS_VTL_pv W=0.090000U L='LMIN_pv'
M_i_32 GNDx RN net_005 GNDx NMOS_VTL_pv W=0.090000U L='LMIN_pv'
M_i_38 GNDx net_003 net_006 GNDx NMOS_VTL_pv W=0.210000U L='LMIN_pv'
M_i_45 net_007 net_003 GNDx GNDx NMOS_VTL_pv W=0.210000U L='LMIN_pv'
M_i_49 net_008 net_001 net_007 GNDx NMOS_VTL_pv W=0.210000U L='LMIN_pv'
M_i_55 net_009 net_000 net_008 GNDx NMOS_VTL_pv W=0.090000U L='LMIN_pv'
M_i_59 GNDx net_011 net_009 GNDx NMOS_VTL_pv W=0.090000U L='LMIN_pv'
M_i_65 net_010 RN GNDx GNDx NMOS_VTL_pv W=0.210000U L='LMIN_pv'
M_i_70 net_011 net_008 net_010 GNDx NMOS_VTL_pv W=0.210000U L='LMIN_pv'
M_i_76 GNDx net_008 QN GNDx NMOS_VTL_pv W=0.415000U L='LMIN_pv'
M_i_83 Q net_011 GNDx GNDx NMOS_VTL_pv W=0.415000U L='LMIN_pv'
M_i_89 VDDx CK net_000 VDDx PMOS_VTL_pv W=0.315000U L='LMIN_pv'
M_i_96 net_001 net_000 VDDx VDDx PMOS_VTL_pv W=0.315000U L='LMIN_pv'
M_i_103 net_012 D VDDx VDDx PMOS_VTL_pv W=0.420000U L='LMIN_pv'
M_i_108 net_003 net_001 net_012 VDDx PMOS_VTL_pv W=0.420000U L='LMIN_pv'
M_i_114 net_013 net_000 net_003 VDDx PMOS_VTL_pv W=0.090000U L='LMIN_pv'
M_i_119 VDDx net_006 net_013 VDDx PMOS_VTL_pv W=0.090000U L='LMIN_pv'
M_i_125 net_013 RN VDDx VDDx PMOS_VTL_pv W=0.090000U L='LMIN_pv'
M_i_136 VDDx net_003 net_006 VDDx PMOS_VTL_pv W=0.315000U L='LMIN_pv'
M_i_143 net_015 net_003 VDDx VDDx PMOS_VTL_pv W=0.315000U L='LMIN_pv'
M_i_147 net_008 net_000 net_015 VDDx PMOS_VTL_pv W=0.315000U L='LMIN_pv'
M_i_153 net_016 net_001 net_008 VDDx PMOS_VTL_pv W=0.090000U L='LMIN_pv'
M_i_159 VDDx net_011 net_016 VDDx PMOS_VTL_pv W=0.090000U L='LMIN_pv'
M_i_165 net_011 RN VDDx VDDx PMOS_VTL_pv W=0.315000U L='LMIN_pv'
M_i_172 VDDx net_008 net_011 VDDx PMOS_VTL_pv W=0.315000U L='LMIN_pv'
M_i_180 VDDx net_008 QN VDDx PMOS_VTL_pv W=0.630000U L='LMIN_pv'
M_i_187 Q net_011 VDDx VDDx PMOS_VTL_pv W=0.630000U L='LMIN_pv'
.ENDS 

**Ringoscillator
XNand1 reset io21 io1 VDD GND NAND2_X1

Xinv2 io1 io2 VDD GND INV_X1
Xinv3 io2 io3 VDD GND INV_X1
Xinv4 io3 io4 VDD GND INV_X1
Xinv5 io4 io5 VDD GND INV_X1
Xinv6 io5 io6 VDD GND INV_X1
Xinv7 io6 io7 VDD GND INV_X1
Xinv8 io7 io8 VDD GND INV_X1
Xinv9 io8 io9 VDD GND INV_X1
Xinv10 io9 io10 VDD GND INV_X1
Xinv11 io10 io11 VDD GND INV_X1
Xinv12 io11 io12 VDD GND INV_X1
Xinv13 io12 io13 VDD GND INV_X1
Xinv14 io13 io14 VDD GND INV_X1
Xinv15 io14 io15 VDD GND INV_X1
Xinv16 io15 io16 VDD GND INV_X1
Xinv17 io16 io17 VDD GND INV_X1
Xinv18 io17 io18 VDD GND INV_X1
Xinv19 io18 io19 VDD GND INV_X1
Xinv20 io19 io20 VDD GND INV_X1
Xinv21 io20 io21 VDD GND INV_X1

**Counter

XDFF0 QN0 io21 reset Q0 QN0 VDD GND DFFR_X1
XDFF1 QN1 QN0 reset Q1 QN1 VDD GND DFFR_X1
XDFF2 QN2 QN1 reset Q2 QN2 VDD GND DFFR_X1
XDFF3 QN3 QN2 reset Q3 QN3 VDD GND DFFR_X1
XDFF4 QN4 QN3 reset Q4 QN4 VDD GND DFFR_X1
XDFF5 QN5 QN4 reset Q5 QN5 VDD GND DFFR_X1
XDFF6 QN6 QN5 reset Q6 QN6 VDD GND DFFR_X1
XDFF7 QN7 QN6 reset Q7 QN7 VDD GND DFFR_X1
XDFF8 QN8 QN7 reset Q8 QN8 VDD GND DFFR_X1
XDFF9 QN9 QN8 reset Q9 QN9 VDD GND DFFR_X1

**register  
XRDFF0 Q0 CLK reset QR0 QRN0 VDD GND DFFR_X1
XRDFF1 Q1 CLK reset QR1 QRN1 VDD GND DFFR_X1
XRDFF2 Q2 CLK reset QR2 QRN2 VDD GND DFFR_X1
XRDFF3 Q3 CLK reset QR3 QRN3 VDD GND DFFR_X1
XRDFF4 Q4 CLK reset QR4 QRN4 VDD GND DFFR_X1
XRDFF5 Q5 CLK reset QR5 QRN5 VDD GND DFFR_X1
XRDFF6 Q6 CLK reset QR6 QRN6 VDD GND DFFR_X1
XRDFF7 Q7 CLK reset QR7 QRN7 VDD GND DFFR_X1
XRDFF8 Q8 CLK reset QR8 QRN8 VDD GND DFFR_X1
XRDFF9 Q9 CLK reset QR9 QRN9 VDD GND DFFR_X1  


* The monitoring
.PRINT TRAN V(QR0) V(QR1) V(QR2) V(QR3) V(QR4) V(QR5) V(QR6) V(QR7) V(QR8) V(QR9)



.END