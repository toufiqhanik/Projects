`timescale 1ns / 1ps

module aes_top(clk,encodedtext);
    input clk;
    output [127:0] encodedtext;
	 
	 wire [127:0] encodedtext;

wire [127:0] tempout;

//clk, plaintextin, keyin, cipertex

aes1 aesencd (.clk(clk),.plaintextin(128'h 54776F204F6E65204E696E652054776F),.keyin(128'h 5468617473206D79204B756E67204675),.cipertex(tempout));

//aes aesencd(.clk(clk),.plaintextin(128'b 01010100011101110110111100100000010011110110111001100101001000000100111001101001011011100110010100100000010101000111011101101111),.keyin(128'b 01010100011010000110000101110100011100110010000001101101011110010010000001001011011101010110111001100111001000000100011001110101),.cipertex(tempout));

assign encodedtext = tempout[127:0];

endmodule
