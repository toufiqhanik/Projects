.Option ingold=2 accurate
.OPTION MEASDGT=8
.OPTION NUMDGT=10
+ RUNLVL=5 ACCURATE
.op
.PARAM LMIN='50E-9'
.PARAM VDD_VALUE=1.2
.PARAM VDD_HALF=0.6
.OPTION BRIEF=1

.OPTION POST=2
.OPTION MEASFORM=3
.OPTION PROBE=1

VSUPPLY VDD 0 VDD_VALUE
VSUPPLYGND GND 0 0
.TRAN 10p 7N START=0N

.include './trans_model_nk'
.temp 25

X0 A0    N3 VDD GND INV_X1
X1 A2 A1 T1 VDD GND XOR2_X1
X2 A2 T1 T2 VDD GND AND2_x1
X3 A3 T2 T3 VDD GND XOR2_X1
X4 A0 T3 Y0 VDD GND XOR2_X1
X5 T1 T3 T4 VDD GND AND2_X1
X6 T1 Y0 T5 VDD GND XOR2_X1
X7 T4 A2 T6 VDD GND XOR2_X1
X8 A0 T6 T7 VDD GND OR2_X1
X9 T5 T7 Y1 VDD GND XOR2_X1
XA T6 N3 T8 VDD GND XOR2_X1
XB Y1 T8 Y3 VDD GND XOR2_X1
XC T5 T8 T9 VDD GND OR2_X1
XD T3 T9 Y2 VDD GND XOR2_X1

***add round key
*.PARAM ki3 = 0
*.PARAM ki2 = 0
*.PARAM ki1 = 0
*.PARAM ki0 = VDD_VALUE


Xxor3 Ak3 VDD_VALUE A3 VDD GND XOR2_X1
Xxor2 Ak2 VDD_VALUE A2 VDD GND XOR2_X1
Xxor1 Ak1 VDD_VALUE A1 VDD GND XOR2_X1
Xxor0 Ak0 0 A0 VDD GND XOR2_X1




***registers

Vinputclk CLK GND PWL (0 0 4.999n 0 5n VDD_VALUE 7n VDD_VALUE)

**Vinputrst reset GND PWL(0 VDD_VALUE 0.2n VDD_VALUE 0.3n 0 1.3n 0 1.4n VDD_VALUE)
Vinputrst reset GND PWL(0 0 1.999n 0 2n VDD_VALUE)  
**falling edge reset


XRDFF0 Y0 CLK reset QR0 QRN0 VDD GND DFFR_X1
XRDFF1 Y1 CLK reset QR1 QRN1 VDD GND DFFR_X1
XRDFF2 Y2 CLK reset QR2 QRN2 VDD GND DFFR_X1
XRDFF3 Y3 CLK reset QR3 QRN3 VDD GND DFFR_X1



*******


*****************************
* The subcircuit for AND
.SUBCKT AND2_X1
+ A1 A2
+ ZN
+ VDD GND
M_i_2 net_0 A2 ZN_neg GND NMOS_VTL W=0.210000U L='LMIN'
M_i_3 GND A1 net_0 GND NMOS_VTL W=0.210000U L='LMIN'
M_i_0 ZN ZN_neg GND GND NMOS_VTL W=0.415000U L='LMIN'
M_i_10 ZN_neg A1 VDD VDD PMOS_VTL W=0.315000U L='LMIN'
M_i_11 VDD A2 ZN_neg VDD PMOS_VTL W=0.315000U L='LMIN'
M_i_1 ZN ZN_neg VDD VDD PMOS_VTL W=0.630000U L='LMIN'
.ENDS


******** OR MODEL ***********
* The subcircuit for OR
.SUBCKT OR2_X1
+ A1 A2
+ ZN
+ VDD GND
M_i_2 ZN_neg A1 GND GND NMOS_VTL W=0.210000U L='LMIN'
M_i_3 GND A2 ZN_neg GND NMOS_VTL W=0.210000U L='LMIN'
M_i_0 ZN ZN_neg GND GND NMOS_VTL W=0.415000U L='LMIN'
M_i_10 net_0 A1 ZN_neg VDD PMOS_VTL W=0.315000U L='LMIN'
M_i_11 VDD A2 net_0 VDD PMOS_VTL W=0.315000U L='LMIN'
M_i_1 ZN ZN_neg VDD VDD PMOS_VTL W=0.630000U L='LMIN'
.ENDS

******** INV MODEL ***********
* The subcircuit for INV
.SUBCKT INV_X1
+ A
+ ZN
+ VDD GND
M_i_0 ZN A GND GND NMOS_VTL W=0.415000U L='LMIN'
M_i_10 ZN A VDD VDD PMOS_VTL W=0.630000U L='LMIN'
.ENDS

******** XOR MODEL ***********
* The subcircuit for XOR
.SUBCKT XOR2_X1
+ A B
+ Z
+ VDD GND
M_i_0 net_000 A GND GND NMOS_VTL W=0.210000U L='LMIN'
M_i_7 GND B net_000 GND NMOS_VTL W=0.210000U L='LMIN'
M_i_13 Z net_000 GND GND NMOS_VTL W=0.415000U L='LMIN'
M_i_19 net_001 A Z GND NMOS_VTL W=0.415000U L='LMIN'
M_i_24 GND B net_001 GND NMOS_VTL W=0.415000U L='LMIN'
M_i_10 net_002 A net_000 VDD PMOS_VTL W=0.315000U L='LMIN'
M_i_11 VDD B net_002 VDD PMOS_VTL W=0.315000U L='LMIN'
M_i_41 net_003 net_000 VDD VDD PMOS_VTL W=0.630000U L='LMIN'
M_i_20 Z A net_003 VDD PMOS_VTL W=0.630000U L='LMIN'
M_i_21 net_003 B Z VDD PMOS_VTL W=0.630000U L='LMIN'

.ENDS
****************************

******** DFFR_X1 MODEL ***********
* The subcircuit for DFFR_X1
.SUBCKT DFFR_X1
+ D CK RN
+ Q QN
+ VDDx GNDx

*.PININFO D:I RN:I CK:I Q:O QN:O VDDx:P GNDx:G 
M_i_0 GNDx CK net_000 GNDx NMOS_VTL W=0.210000U L='LMIN'
M_i_7 net_001 net_000 GNDx GNDx NMOS_VTL W=0.210000U L='LMIN'
M_i_13 net_002 D GNDx GNDx NMOS_VTL W=0.275000U L='LMIN'
M_i_18 net_003 net_000 net_002 GNDx NMOS_VTL W=0.275000U L='LMIN'
M_i_24 net_004 net_001 net_003 GNDx NMOS_VTL W=0.090000U L='LMIN'
M_i_28 net_005 net_006 net_004 GNDx NMOS_VTL W=0.090000U L='LMIN'
M_i_32 GNDx RN net_005 GNDx NMOS_VTL W=0.090000U L='LMIN'
M_i_38 GNDx net_003 net_006 GNDx NMOS_VTL W=0.210000U L='LMIN'
M_i_45 net_007 net_003 GNDx GNDx NMOS_VTL W=0.210000U L='LMIN'
M_i_49 net_008 net_001 net_007 GNDx NMOS_VTL W=0.210000U L='LMIN'
M_i_55 net_009 net_000 net_008 GNDx NMOS_VTL W=0.090000U L='LMIN'
M_i_59 GNDx net_011 net_009 GNDx NMOS_VTL W=0.090000U L='LMIN'
M_i_65 net_010 RN GNDx GNDx NMOS_VTL W=0.210000U L='LMIN'
M_i_70 net_011 net_008 net_010 GNDx NMOS_VTL W=0.210000U L='LMIN'
M_i_76 GNDx net_008 QN GNDx NMOS_VTL W=0.415000U L='LMIN'
M_i_83 Q net_011 GNDx GNDx NMOS_VTL W=0.415000U L='LMIN'
M_i_89 VDDx CK net_000 VDDx PMOS_VTL W=0.315000U L='LMIN'
M_i_96 net_001 net_000 VDDx VDDx PMOS_VTL W=0.315000U L='LMIN'
M_i_103 net_012 D VDDx VDDx PMOS_VTL W=0.420000U L='LMIN'
M_i_108 net_003 net_001 net_012 VDDx PMOS_VTL W=0.420000U L='LMIN'
M_i_114 net_013 net_000 net_003 VDDx PMOS_VTL W=0.090000U L='LMIN'
M_i_119 VDDx net_006 net_013 VDDx PMOS_VTL W=0.090000U L='LMIN'
M_i_125 net_013 RN VDDx VDDx PMOS_VTL W=0.090000U L='LMIN'
M_i_136 VDDx net_003 net_006 VDDx PMOS_VTL W=0.315000U L='LMIN'
M_i_143 net_015 net_003 VDDx VDDx PMOS_VTL W=0.315000U L='LMIN'
M_i_147 net_008 net_000 net_015 VDDx PMOS_VTL W=0.315000U L='LMIN'
M_i_153 net_016 net_001 net_008 VDDx PMOS_VTL W=0.090000U L='LMIN'
M_i_159 VDDx net_011 net_016 VDDx PMOS_VTL W=0.090000U L='LMIN'
M_i_165 net_011 RN VDDx VDDx PMOS_VTL W=0.315000U L='LMIN'
M_i_172 VDDx net_008 net_011 VDDx PMOS_VTL W=0.315000U L='LMIN'
M_i_180 VDDx net_008 QN VDDx PMOS_VTL W=0.630000U L='LMIN'
M_i_187 Q net_011 VDDx VDDx PMOS_VTL W=0.630000U L='LMIN'
.ENDS 
***********************

.PARAM A3i = 0
.PARAM A2i = 0
.PARAM A1i = 0
.PARAM A0i = 0


VA3 Ak3 0 PWL (0ns 0 2.499ns 0 2.5ns A3i 7ns A3i)
VA2 Ak2 0 PWL (0ns 0 2.499ns 0 2.5ns A2i 7ns A2i)
VA1 Ak1 0 PWL (0ns 0 2.499ns 0 2.5ns A1i 7ns A1i)
VA0 Ak0 0 PWL (0ns 0 2.499ns 0 2.5ns A0i 7ns A0i)

* The monitoring
.PROBE TRAN V(A0) V(A1) V(A2) V(A3) V(Y0) V(Y1) V(Y2) V(Y3) V(QR0) V(QR1) V(QR2) V(QR3) V(reset) V(CLK) V(Ak0) V(Ak1) V(Ak2) V(Ak3) 
.PRINT TRAN V(A0) V(A1) V(A2) V(A3) V(Y0) V(Y1) V(Y2) V(Y3) V(QR0) V(QR1) V(QR2) V(QR3) V(reset) V(CLK) V(Ak0) V(Ak1) V(Ak2) V(Ak3) 
.PRINT Pvdd=PAR('-VDD_VALUE*I(VSUPPLY)')
.PROBE Pvdd=PAR('-VDD_VALUE*I(VSUPPLY)')


.ALTER
.PARAM A3i=0 A2i=0 A1i=0 A0i=VDD_VALUE 

.ALTER
.PARAM A3i=0 A2i=0 A1i=VDD_VALUE A0i=0 

.ALTER
.PARAM A3i=0 A2i=0 A1i=VDD_VALUE A0i=VDD_VALUE 

.ALTER
.PARAM A3i=0 A2i=VDD_VALUE A1i=0 A0i=0 

.ALTER
.PARAM A3i=0 A2i=VDD_VALUE A1i=0 A0i=VDD_VALUE 

.ALTER
.PARAM A3i=0 A2i=VDD_VALUE A1i=VDD_VALUE A0i=0 

.ALTER
.PARAM A3i=0 A2i=VDD_VALUE A1i=VDD_VALUE A0i=VDD_VALUE 

.ALTER
.PARAM A3i=VDD_VALUE A2i=0 A1i=0 A0i=0 

.ALTER
.PARAM A3i=VDD_VALUE A2i=0 A1i=0 A0i=VDD_VALUE 

.ALTER
.PARAM A3i=VDD_VALUE A2i=0 A1i=VDD_VALUE A0i=0 

.ALTER
.PARAM A3i=VDD_VALUE A2i=0 A1i=VDD_VALUE A0i=VDD_VALUE 

.ALTER
.PARAM A3i=VDD_VALUE A2i=VDD_VALUE A1i=0 A0i=0 

.ALTER
.PARAM A3i=VDD_VALUE A2i=VDD_VALUE A1i=0 A0i=VDD_VALUE 

.ALTER
.PARAM A3i=VDD_VALUE A2i=VDD_VALUE A1i=VDD_VALUE A0i=0 

.ALTER
.PARAM A3i=VDD_VALUE A2i=VDD_VALUE A1i=VDD_VALUE A0i=VDD_VALUE 

.END