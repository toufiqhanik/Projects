module c1908 (N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,N94,N99,N104,N2753,N2754,N2755,N2756,N2762,N2767,N2768,N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2811,N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2899);
input N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,N94,N99,N104;
output N2753,N2754,N2755,N2756,N2762,N2767,N2768,N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2811,N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2899;
wire N190,N194,N197,N201,N206,N209,N212,N216,N220,N225,N229,N232,N235,N239,N243,N247,N251,N252,N253,N256,N257,N260,N263,N266,N269,N272,N275,N276,N277,N280,N283,N290,N297,N300,N303,N306,N313,N316,N319,N326,N331,N338,N343,N346,N349,N352,N355,N358,N361,N364,N367,N370,N373,N376,N379,N382,N385,N388,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N559,N562,N565,N568,N571,N574,N577,N580,N583,N586,N589,N592,N595,N598,N601,N602,N603,N608,N612,N616,N619,N622,N625,N628,N631,N634,N637,N640,N643,N646,N649,N652,N655,N658,N661,N664,N667,N670,N673,N676,N679,N682,N685,N688,N691,N694,N697,N700,N703,N706,N709,N712,N715,N718,N721,N724,N727,N730,N733,N736,N739,N742,N745,N748,N751,N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,N903,N907,N910,N913,N914,N915,N916,N917,N918,N919,N920,N921,N922,N923,N926,N935,N938,N939,N942,N943,N946,N947,N950,N951,N954,N955,N958,N959,N962,N965,N968,N969,N972,N973,N976,N977,N980,N981,N984,N985,N988,N989,N990,N991,N992,N993,N994,N997,N998,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1013,N1016,N1019,N1022,N1025,N1028,N1031,N1034,N1037,N1040,N1043,N1046,N1049,N1054,N1055,N1063,N1064,N1067,N1068,N1119,N1120,N1121,N1122,N1128,N1129,N1130,N1131,N1132,N1133,N1148,N1149,N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1167,N1168,N1171,N1188,N1205,N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1235,N1238,N1239,N1240,N1241,N1242,N1243,N1246,N1249,N1252,N1255,N1258,N1261,N1264,N1267,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,N1317,N1318,N1319,N1322,N1327,N1328,N1334,N1344,N1345,N1346,N1348,N1349,N1350,N1351,N1352,N1355,N1358,N1361,N1364,N1367,N1370,N1373,N1376,N1379,N1383,N1386,N1387,N1388,N1389,N1390,N1393,N1396,N1397,N1398,N1399,N1409,N1412,N1413,N1416,N1419,N1433,N1434,N1438,N1439,N1440,N1443,N1444,N1445,N1446,N1447,N1448,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,N1463,N1464,N1468,N1469,N1470,N1471,N1472,N1475,N1476,N1478,N1481,N1484,N1487,N1488,N1489,N1490,N1491,N1492,N1493,N1494,N1495,N1496,N1498,N1499,N1500,N1501,N1504,N1510,N1513,N1514,N1517,N1520,N1521,N1522,N1526,N1527,N1528,N1529,N1530,N1531,N1532,N1534,N1537,N1540,N1546,N1554,N1557,N1561,N1567,N1568,N1569,N1571,N1576,N1588,N1591,N1593,N1594,N1595,N1596,N1600,N1603,N1606,N1609,N1612,N1615,N1620,N1623,N1635,N1636,N1638,N1639,N1640,N1643,N1647,N1651,N1658,N1661,N1664,N1671,N1672,N1675,N1677,N1678,N1679,N1680,N1681,N1682,N1683,N1685,N1688,N1697,N1701,N1706,N1707,N1708,N1709,N1710,N1711,N1712,N1713,N1714,N1717,N1720,N1721,N1723,N1727,N1728,N1730,N1731,N1734,N1740,N1741,N1742,N1746,N1747,N1748,N1751,N1759,N1761,N1762,N1763,N1764,N1768,N1769,N1772,N1773,N1774,N1777,N1783,N1784,N1785,N1786,N1787,N1788,N1791,N1792,N1795,N1796,N1798,N1801,N1802,N1807,N1808,N1809,N1810,N1812,N1815,N1818,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1830,N1837,N1838,N1841,N1848,N1849,N1850,N1852,N1855,N1856,N1857,N1858,N1864,N1865,N1866,N1869,N1872,N1875,N1878,N1879,N1882,N1883,N1884,N1885,N1889,N1895,N1896,N1897,N1898,N1902,N1910,N1911,N1912,N1913,N1915,N1919,N1920,N1921,N1922,N1923,N1924,N1927,N1930,N1933,N1936,N1937,N1938,N1941,N1942,N1944,N1947,N1950,N1953,N1958,N1961,N1965,N1968,N1975,N1976,N1977,N1978,N1979,N1980,N1985,N1987,N1999,N2000,N2002,N2003,N2004,N2005,N2006,N2007,N2008,N2009,N2012,N2013,N2014,N2015,N2016,N2018,N2019,N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2030,N2033,N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2047,N2052,N2055,N2060,N2061,N2062,N2067,N2068,N2071,N2076,N2077,N2078,N2081,N2086,N2089,N2104,N2119,N2129,N2143,N2148,N2151,N2196,N2199,N2202,N2205,N2214,N2215,N2216,N2217,N2222,N2223,N2224,N2225,N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,N2236,N2237,N2240,N2241,N2244,N2245,N2250,N2253,N2256,N2257,N2260,N2263,N2266,N2269,N2272,N2279,N2286,N2297,N2315,N2326,N2340,N2353,N2361,N2375,N2384,N2385,N2386,N2426,N2427,N2537,N2540,N2543,N2546,N2549,N2552,N2555,N2558,N2561,N2564,N2567,N2570,N2573,N2576,N2594,N2597,N2600,N2603,N2606,N2611,N2614,N2617,N2620,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,N2639,N2642,N2645,N2648,N2651,N2655,N2658,N2661,N2664,N2669,N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2682,N2683,N2688,N2689,N2690,N2691,N2710,N2720,N2721,N2722,N2723,N2724,N2725,N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,N2746,N2747,N2750,N2757,N2758,N2759,N2760,N2761,N2763,N2764,N2765,N2766,N2773,N2776,N2788,N2789,N2800,N2807,N2808,N2809,N2810,N2812,N2815,N2818,N2821,N2824,N2827,N2828,N2829,N2843,N2846,N2850,N2851,N2852,N2853,N2854,N2857,N2858,N2859,N2860,N2861,N2862,N2863,N2866,N2867,N2868,N2869,N2870,N2871,N2872,N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,N2883,N2895,N2896,N2897,N2898;
INVX1 NOT1_1 (.Y(N190),.A(N1));
INVX1 NOT1_2 (.Y(N194),.A(N4));
INVX1 NOT1_3 (.Y(N197),.A(N7));
INVX1 NOT1_4 (.Y(N201),.A(N10));
INVX1 NOT1_5 (.Y(N206),.A(N13));
INVX1 NOT1_6 (.Y(N209),.A(N16));
INVX1 NOT1_7 (.Y(N212),.A(N19));
INVX1 NOT1_8 (.Y(N216),.A(N22));
INVX1 NOT1_9 (.Y(N220),.A(N25));
INVX1 NOT1_10 (.Y(N225),.A(N28));
INVX1 NOT1_11 (.Y(N229),.A(N31));
INVX1 NOT1_12 (.Y(N232),.A(N34));
INVX1 NOT1_13 (.Y(N235),.A(N37));
INVX1 NOT1_14 (.Y(N239),.A(N40));
INVX1 NOT1_15 (.Y(N243),.A(N43));
INVX1 NOT1_16 (.Y(N247),.A(N46));
NAND2X1 NAND2_17 (.Y(N251),.A(N63),.B(N88));
NAND2X1 NAND2_18 (.Y(N252),.A(N66),.B(N91));
INVX1 NOT1_19 (.Y(N253),.A(N72));
INVX1 NOT1_20 (.Y(N256),.A(N72));
BUFX1 BUFF1_21 (.Y(N257),.A(N69));
BUFX1 BUFF1_22 (.Y(N260),.A(N69));
INVX1 NOT1_23 (.Y(N263),.A(N76));
INVX1 NOT1_24 (.Y(N266),.A(N79));
INVX1 NOT1_25 (.Y(N269),.A(N82));
INVX1 NOT1_26 (.Y(N272),.A(N85));
INVX1 NOT1_27 (.Y(N275),.A(N104));
INVX1 NOT1_28 (.Y(N276),.A(N104));
INVX1 NOT1_29 (.Y(N277),.A(N88));
INVX1 NOT1_30 (.Y(N280),.A(N91));
BUFX1 BUFF1_31 (.Y(N283),.A(N94));
INVX1 NOT1_32 (.Y(N290),.A(N94));
BUFX1 BUFF1_33 (.Y(N297),.A(N94));
INVX1 NOT1_34 (.Y(N300),.A(N94));
BUFX1 BUFF1_35 (.Y(N303),.A(N99));
INVX1 NOT1_36 (.Y(N306),.A(N99));
INVX1 NOT1_37 (.Y(N313),.A(N99));
BUFX1 BUFF1_38 (.Y(N316),.A(N104));
INVX1 NOT1_39 (.Y(N319),.A(N104));
BUFX1 BUFF1_40 (.Y(N326),.A(N104));
BUFX1 BUFF1_41 (.Y(N331),.A(N104));
INVX1 NOT1_42 (.Y(N338),.A(N104));
BUFX1 BUFF1_43 (.Y(N343),.A(N1));
BUFX1 BUFF1_44 (.Y(N346),.A(N4));
BUFX1 BUFF1_45 (.Y(N349),.A(N7));
BUFX1 BUFF1_46 (.Y(N352),.A(N10));
BUFX1 BUFF1_47 (.Y(N355),.A(N13));
BUFX1 BUFF1_48 (.Y(N358),.A(N16));
BUFX1 BUFF1_49 (.Y(N361),.A(N19));
BUFX1 BUFF1_50 (.Y(N364),.A(N22));
BUFX1 BUFF1_51 (.Y(N367),.A(N25));
BUFX1 BUFF1_52 (.Y(N370),.A(N28));
BUFX1 BUFF1_53 (.Y(N373),.A(N31));
BUFX1 BUFF1_54 (.Y(N376),.A(N34));
BUFX1 BUFF1_55 (.Y(N379),.A(N37));
BUFX1 BUFF1_56 (.Y(N382),.A(N40));
BUFX1 BUFF1_57 (.Y(N385),.A(N43));
BUFX1 BUFF1_58 (.Y(N388),.A(N46));
INVX1 NOT1_59 (.Y(N534),.A(N343));
INVX1 NOT1_60 (.Y(N535),.A(N346));
INVX1 NOT1_61 (.Y(N536),.A(N349));
INVX1 NOT1_62 (.Y(N537),.A(N352));
INVX1 NOT1_63 (.Y(N538),.A(N355));
INVX1 NOT1_64 (.Y(N539),.A(N358));
INVX1 NOT1_65 (.Y(N540),.A(N361));
INVX1 NOT1_66 (.Y(N541),.A(N364));
INVX1 NOT1_67 (.Y(N542),.A(N367));
INVX1 NOT1_68 (.Y(N543),.A(N370));
INVX1 NOT1_69 (.Y(N544),.A(N373));
INVX1 NOT1_70 (.Y(N545),.A(N376));
INVX1 NOT1_71 (.Y(N546),.A(N379));
INVX1 NOT1_72 (.Y(N547),.A(N382));
INVX1 NOT1_73 (.Y(N548),.A(N385));
INVX1 NOT1_74 (.Y(N549),.A(N388));
NAND2X1 NAND2_75 (.Y(N550),.A(N306),.B(N331));
NAND2X1 NAND2_76 (.Y(N551),.A(N306),.B(N331));
NAND2X1 NAND2_77 (.Y(N552),.A(N306),.B(N331));
NAND2X1 NAND2_78 (.Y(N553),.A(N306),.B(N331));
NAND2X1 NAND2_79 (.Y(N554),.A(N306),.B(N331));
NAND2X1 NAND2_80 (.Y(N555),.A(N306),.B(N331));
BUFX1 BUFF1_81 (.Y(N556),.A(N190));
BUFX1 BUFF1_82 (.Y(N559),.A(N194));
BUFX1 BUFF1_83 (.Y(N562),.A(N206));
BUFX1 BUFF1_84 (.Y(N565),.A(N209));
BUFX1 BUFF1_85 (.Y(N568),.A(N225));
BUFX1 BUFF1_86 (.Y(N571),.A(N243));
AND2X1 AND2_87 (.Y(N574),.A(N63),.B(N319));
BUFX1 BUFF1_88 (.Y(N577),.A(N220));
BUFX1 BUFF1_89 (.Y(N580),.A(N229));
BUFX1 BUFF1_90 (.Y(N583),.A(N232));
AND2X1 AND2_91 (.Y(N586),.A(N66),.B(N319));
BUFX1 BUFF1_92 (.Y(N589),.A(N239));
AND2X1 AND_tmp1 (.Y(ttmp1),.A(N253),.B(N319));
AND2X1 AND_tmp2 (.Y(N592),.A(N49),.B(ttmp1));
BUFX1 BUFF1_94 (.Y(N595),.A(N247));
BUFX1 BUFF1_95 (.Y(N598),.A(N239));
NAND2X1 NAND2_96 (.Y(N601),.A(N326),.B(N277));
NAND2X1 NAND2_97 (.Y(N602),.A(N326),.B(N280));
NAND2X1 NAND2_98 (.Y(N603),.A(N260),.B(N72));
NAND2X1 NAND2_99 (.Y(N608),.A(N260),.B(N300));
NAND2X1 NAND2_100 (.Y(N612),.A(N256),.B(N300));
BUFX1 BUFF1_101 (.Y(N616),.A(N201));
BUFX1 BUFF1_102 (.Y(N619),.A(N216));
BUFX1 BUFF1_103 (.Y(N622),.A(N220));
BUFX1 BUFF1_104 (.Y(N625),.A(N239));
BUFX1 BUFF1_105 (.Y(N628),.A(N190));
BUFX1 BUFF1_106 (.Y(N631),.A(N190));
BUFX1 BUFF1_107 (.Y(N634),.A(N194));
BUFX1 BUFF1_108 (.Y(N637),.A(N229));
BUFX1 BUFF1_109 (.Y(N640),.A(N197));
AND2X1 AND_tmp3 (.Y(ttmp3),.A(N257),.B(N319));
AND2X1 AND_tmp4 (.Y(N643),.A(N56),.B(ttmp3));
BUFX1 BUFF1_111 (.Y(N646),.A(N232));
BUFX1 BUFF1_112 (.Y(N649),.A(N201));
BUFX1 BUFF1_113 (.Y(N652),.A(N235));
AND2X1 AND_tmp5 (.Y(ttmp5),.A(N257),.B(N319));
AND2X1 AND_tmp6 (.Y(N655),.A(N60),.B(ttmp5));
BUFX1 BUFF1_115 (.Y(N658),.A(N263));
BUFX1 BUFF1_116 (.Y(N661),.A(N263));
BUFX1 BUFF1_117 (.Y(N664),.A(N266));
BUFX1 BUFF1_118 (.Y(N667),.A(N266));
BUFX1 BUFF1_119 (.Y(N670),.A(N269));
BUFX1 BUFF1_120 (.Y(N673),.A(N269));
BUFX1 BUFF1_121 (.Y(N676),.A(N272));
BUFX1 BUFF1_122 (.Y(N679),.A(N272));
AND2X1 AND2_123 (.Y(N682),.A(N251),.B(N316));
AND2X1 AND2_124 (.Y(N685),.A(N252),.B(N316));
BUFX1 BUFF1_125 (.Y(N688),.A(N197));
BUFX1 BUFF1_126 (.Y(N691),.A(N197));
BUFX1 BUFF1_127 (.Y(N694),.A(N212));
BUFX1 BUFF1_128 (.Y(N697),.A(N212));
BUFX1 BUFF1_129 (.Y(N700),.A(N247));
BUFX1 BUFF1_130 (.Y(N703),.A(N247));
BUFX1 BUFF1_131 (.Y(N706),.A(N235));
BUFX1 BUFF1_132 (.Y(N709),.A(N235));
BUFX1 BUFF1_133 (.Y(N712),.A(N201));
BUFX1 BUFF1_134 (.Y(N715),.A(N201));
BUFX1 BUFF1_135 (.Y(N718),.A(N206));
BUFX1 BUFF1_136 (.Y(N721),.A(N216));
AND2X1 AND_tmp7 (.Y(ttmp7),.A(N253),.B(N319));
AND2X1 AND_tmp8 (.Y(N724),.A(N53),.B(ttmp7));
BUFX1 BUFF1_138 (.Y(N727),.A(N243));
BUFX1 BUFF1_139 (.Y(N730),.A(N220));
BUFX1 BUFF1_140 (.Y(N733),.A(N220));
BUFX1 BUFF1_141 (.Y(N736),.A(N209));
BUFX1 BUFF1_142 (.Y(N739),.A(N216));
BUFX1 BUFF1_143 (.Y(N742),.A(N225));
BUFX1 BUFF1_144 (.Y(N745),.A(N243));
BUFX1 BUFF1_145 (.Y(N748),.A(N212));
BUFX1 BUFF1_146 (.Y(N751),.A(N225));
INVX1 NOT1_147 (.Y(N886),.A(N682));
INVX1 NOT1_148 (.Y(N887),.A(N685));
INVX1 NOT1_149 (.Y(N888),.A(N616));
INVX1 NOT1_150 (.Y(N889),.A(N619));
INVX1 NOT1_151 (.Y(N890),.A(N622));
INVX1 NOT1_152 (.Y(N891),.A(N625));
INVX1 NOT1_153 (.Y(N892),.A(N631));
INVX1 NOT1_154 (.Y(N893),.A(N643));
INVX1 NOT1_155 (.Y(N894),.A(N649));
INVX1 NOT1_156 (.Y(N895),.A(N652));
INVX1 NOT1_157 (.Y(N896),.A(N655));
AND2X1 AND2_158 (.Y(N897),.A(N49),.B(N612));
AND2X1 AND2_159 (.Y(N898),.A(N56),.B(N608));
NAND2X1 NAND2_160 (.Y(N899),.A(N53),.B(N612));
NAND2X1 NAND2_161 (.Y(N903),.A(N60),.B(N608));
NAND2X1 NAND2_162 (.Y(N907),.A(N49),.B(N612));
NAND2X1 NAND2_163 (.Y(N910),.A(N56),.B(N608));
INVX1 NOT1_164 (.Y(N913),.A(N661));
INVX1 NOT1_165 (.Y(N914),.A(N658));
INVX1 NOT1_166 (.Y(N915),.A(N667));
INVX1 NOT1_167 (.Y(N916),.A(N664));
INVX1 NOT1_168 (.Y(N917),.A(N673));
INVX1 NOT1_169 (.Y(N918),.A(N670));
INVX1 NOT1_170 (.Y(N919),.A(N679));
INVX1 NOT1_171 (.Y(N920),.A(N676));
AND2X1 AND_tmp9 (.Y(ttmp9),.A(N326),.B(N603));
AND2X1 AND_tmp10 (.Y(ttmp10),.A(N277),.B(ttmp9));
NAND2X1 NAND_tmp11 (.Y(N921),.A(N297),.B(ttmp10));
AND2X1 AND_tmp12 (.Y(ttmp12),.A(N326),.B(N603));
AND2X1 AND_tmp13 (.Y(ttmp13),.A(N280),.B(ttmp12));
NAND2X1 NAND_tmp14 (.Y(N922),.A(N297),.B(ttmp13));
AND2X1 AND_tmp15 (.Y(ttmp15),.A(N338),.B(N603));
NAND2X1 NAND_tmp16 (.Y(N923),.A(N303),.B(ttmp15));
AND2X1 AND_tmp17 (.Y(ttmp17),.A(N338),.B(N603));
AND2X1 AND_tmp18 (.Y(N926),.A(N303),.B(ttmp17));
BUFX1 BUFF1_176 (.Y(N935),.A(N556));
INVX1 NOT1_177 (.Y(N938),.A(N688));
BUFX1 BUFF1_178 (.Y(N939),.A(N556));
INVX1 NOT1_179 (.Y(N942),.A(N691));
BUFX1 BUFF1_180 (.Y(N943),.A(N562));
INVX1 NOT1_181 (.Y(N946),.A(N694));
BUFX1 BUFF1_182 (.Y(N947),.A(N562));
INVX1 NOT1_183 (.Y(N950),.A(N697));
BUFX1 BUFF1_184 (.Y(N951),.A(N568));
INVX1 NOT1_185 (.Y(N954),.A(N700));
BUFX1 BUFF1_186 (.Y(N955),.A(N568));
INVX1 NOT1_187 (.Y(N958),.A(N703));
BUFX1 BUFF1_188 (.Y(N959),.A(N574));
BUFX1 BUFF1_189 (.Y(N962),.A(N574));
BUFX1 BUFF1_190 (.Y(N965),.A(N580));
INVX1 NOT1_191 (.Y(N968),.A(N706));
BUFX1 BUFF1_192 (.Y(N969),.A(N580));
INVX1 NOT1_193 (.Y(N972),.A(N709));
BUFX1 BUFF1_194 (.Y(N973),.A(N586));
INVX1 NOT1_195 (.Y(N976),.A(N712));
BUFX1 BUFF1_196 (.Y(N977),.A(N586));
INVX1 NOT1_197 (.Y(N980),.A(N715));
BUFX1 BUFF1_198 (.Y(N981),.A(N592));
INVX1 NOT1_199 (.Y(N984),.A(N628));
BUFX1 BUFF1_200 (.Y(N985),.A(N592));
INVX1 NOT1_201 (.Y(N988),.A(N718));
INVX1 NOT1_202 (.Y(N989),.A(N721));
INVX1 NOT1_203 (.Y(N990),.A(N634));
INVX1 NOT1_204 (.Y(N991),.A(N724));
INVX1 NOT1_205 (.Y(N992),.A(N727));
INVX1 NOT1_206 (.Y(N993),.A(N637));
BUFX1 BUFF1_207 (.Y(N994),.A(N595));
INVX1 NOT1_208 (.Y(N997),.A(N730));
BUFX1 BUFF1_209 (.Y(N998),.A(N595));
INVX1 NOT1_210 (.Y(N1001),.A(N733));
INVX1 NOT1_211 (.Y(N1002),.A(N736));
INVX1 NOT1_212 (.Y(N1003),.A(N739));
INVX1 NOT1_213 (.Y(N1004),.A(N640));
INVX1 NOT1_214 (.Y(N1005),.A(N742));
INVX1 NOT1_215 (.Y(N1006),.A(N745));
INVX1 NOT1_216 (.Y(N1007),.A(N646));
INVX1 NOT1_217 (.Y(N1008),.A(N748));
INVX1 NOT1_218 (.Y(N1009),.A(N751));
BUFX1 BUFF1_219 (.Y(N1010),.A(N559));
BUFX1 BUFF1_220 (.Y(N1013),.A(N559));
BUFX1 BUFF1_221 (.Y(N1016),.A(N565));
BUFX1 BUFF1_222 (.Y(N1019),.A(N565));
BUFX1 BUFF1_223 (.Y(N1022),.A(N571));
BUFX1 BUFF1_224 (.Y(N1025),.A(N571));
BUFX1 BUFF1_225 (.Y(N1028),.A(N577));
BUFX1 BUFF1_226 (.Y(N1031),.A(N577));
BUFX1 BUFF1_227 (.Y(N1034),.A(N583));
BUFX1 BUFF1_228 (.Y(N1037),.A(N583));
BUFX1 BUFF1_229 (.Y(N1040),.A(N589));
BUFX1 BUFF1_230 (.Y(N1043),.A(N589));
BUFX1 BUFF1_231 (.Y(N1046),.A(N598));
BUFX1 BUFF1_232 (.Y(N1049),.A(N598));
NAND2X1 NAND2_233 (.Y(N1054),.A(N619),.B(N888));
NAND2X1 NAND2_234 (.Y(N1055),.A(N616),.B(N889));
NAND2X1 NAND2_235 (.Y(N1063),.A(N625),.B(N890));
NAND2X1 NAND2_236 (.Y(N1064),.A(N622),.B(N891));
NAND2X1 NAND2_237 (.Y(N1067),.A(N655),.B(N895));
NAND2X1 NAND2_238 (.Y(N1068),.A(N652),.B(N896));
NAND2X1 NAND2_239 (.Y(N1119),.A(N721),.B(N988));
NAND2X1 NAND2_240 (.Y(N1120),.A(N718),.B(N989));
NAND2X1 NAND2_241 (.Y(N1121),.A(N727),.B(N991));
NAND2X1 NAND2_242 (.Y(N1122),.A(N724),.B(N992));
NAND2X1 NAND2_243 (.Y(N1128),.A(N739),.B(N1002));
NAND2X1 NAND2_244 (.Y(N1129),.A(N736),.B(N1003));
NAND2X1 NAND2_245 (.Y(N1130),.A(N745),.B(N1005));
NAND2X1 NAND2_246 (.Y(N1131),.A(N742),.B(N1006));
NAND2X1 NAND2_247 (.Y(N1132),.A(N751),.B(N1008));
NAND2X1 NAND2_248 (.Y(N1133),.A(N748),.B(N1009));
INVX1 NOT1_249 (.Y(N1148),.A(N939));
INVX1 NOT1_250 (.Y(N1149),.A(N935));
NAND2X1 NAND2_251 (.Y(N1150),.A(N1054),.B(N1055));
INVX1 NOT1_252 (.Y(N1151),.A(N943));
INVX1 NOT1_253 (.Y(N1152),.A(N947));
INVX1 NOT1_254 (.Y(N1153),.A(N955));
INVX1 NOT1_255 (.Y(N1154),.A(N951));
INVX1 NOT1_256 (.Y(N1155),.A(N962));
INVX1 NOT1_257 (.Y(N1156),.A(N969));
INVX1 NOT1_258 (.Y(N1157),.A(N977));
NAND2X1 NAND2_259 (.Y(N1158),.A(N1063),.B(N1064));
INVX1 NOT1_260 (.Y(N1159),.A(N985));
NAND2X1 NAND2_261 (.Y(N1160),.A(N985),.B(N892));
INVX1 NOT1_262 (.Y(N1161),.A(N998));
NAND2X1 NAND2_263 (.Y(N1162),.A(N1067),.B(N1068));
INVX1 NOT1_264 (.Y(N1163),.A(N899));
BUFX1 BUFF1_265 (.Y(N1164),.A(N899));
INVX1 NOT1_266 (.Y(N1167),.A(N903));
BUFX1 BUFF1_267 (.Y(N1168),.A(N903));
NAND2X1 NAND2_268 (.Y(N1171),.A(N921),.B(N923));
NAND2X1 NAND2_269 (.Y(N1188),.A(N922),.B(N923));
INVX1 NOT1_270 (.Y(N1205),.A(N1010));
NAND2X1 NAND2_271 (.Y(N1206),.A(N1010),.B(N938));
INVX1 NOT1_272 (.Y(N1207),.A(N1013));
NAND2X1 NAND2_273 (.Y(N1208),.A(N1013),.B(N942));
INVX1 NOT1_274 (.Y(N1209),.A(N1016));
NAND2X1 NAND2_275 (.Y(N1210),.A(N1016),.B(N946));
INVX1 NOT1_276 (.Y(N1211),.A(N1019));
NAND2X1 NAND2_277 (.Y(N1212),.A(N1019),.B(N950));
INVX1 NOT1_278 (.Y(N1213),.A(N1022));
NAND2X1 NAND2_279 (.Y(N1214),.A(N1022),.B(N954));
INVX1 NOT1_280 (.Y(N1215),.A(N1025));
NAND2X1 NAND2_281 (.Y(N1216),.A(N1025),.B(N958));
INVX1 NOT1_282 (.Y(N1217),.A(N1028));
INVX1 NOT1_283 (.Y(N1218),.A(N959));
INVX1 NOT1_284 (.Y(N1219),.A(N1031));
INVX1 NOT1_285 (.Y(N1220),.A(N1034));
NAND2X1 NAND2_286 (.Y(N1221),.A(N1034),.B(N968));
INVX1 NOT1_287 (.Y(N1222),.A(N965));
INVX1 NOT1_288 (.Y(N1223),.A(N1037));
NAND2X1 NAND2_289 (.Y(N1224),.A(N1037),.B(N972));
INVX1 NOT1_290 (.Y(N1225),.A(N1040));
NAND2X1 NAND2_291 (.Y(N1226),.A(N1040),.B(N976));
INVX1 NOT1_292 (.Y(N1227),.A(N973));
INVX1 NOT1_293 (.Y(N1228),.A(N1043));
NAND2X1 NAND2_294 (.Y(N1229),.A(N1043),.B(N980));
INVX1 NOT1_295 (.Y(N1230),.A(N981));
NAND2X1 NAND2_296 (.Y(N1231),.A(N981),.B(N984));
NAND2X1 NAND2_297 (.Y(N1232),.A(N1119),.B(N1120));
NAND2X1 NAND2_298 (.Y(N1235),.A(N1121),.B(N1122));
INVX1 NOT1_299 (.Y(N1238),.A(N1046));
NAND2X1 NAND2_300 (.Y(N1239),.A(N1046),.B(N997));
INVX1 NOT1_301 (.Y(N1240),.A(N994));
INVX1 NOT1_302 (.Y(N1241),.A(N1049));
NAND2X1 NAND2_303 (.Y(N1242),.A(N1049),.B(N1001));
NAND2X1 NAND2_304 (.Y(N1243),.A(N1128),.B(N1129));
NAND2X1 NAND2_305 (.Y(N1246),.A(N1130),.B(N1131));
NAND2X1 NAND2_306 (.Y(N1249),.A(N1132),.B(N1133));
BUFX1 BUFF1_307 (.Y(N1252),.A(N907));
BUFX1 BUFF1_308 (.Y(N1255),.A(N907));
BUFX1 BUFF1_309 (.Y(N1258),.A(N910));
BUFX1 BUFF1_310 (.Y(N1261),.A(N910));
INVX1 NOT1_311 (.Y(N1264),.A(N1150));
NAND2X1 NAND2_312 (.Y(N1267),.A(N631),.B(N1159));
NAND2X1 NAND2_313 (.Y(N1309),.A(N688),.B(N1205));
NAND2X1 NAND2_314 (.Y(N1310),.A(N691),.B(N1207));
NAND2X1 NAND2_315 (.Y(N1311),.A(N694),.B(N1209));
NAND2X1 NAND2_316 (.Y(N1312),.A(N697),.B(N1211));
NAND2X1 NAND2_317 (.Y(N1313),.A(N700),.B(N1213));
NAND2X1 NAND2_318 (.Y(N1314),.A(N703),.B(N1215));
NAND2X1 NAND2_319 (.Y(N1315),.A(N706),.B(N1220));
NAND2X1 NAND2_320 (.Y(N1316),.A(N709),.B(N1223));
NAND2X1 NAND2_321 (.Y(N1317),.A(N712),.B(N1225));
NAND2X1 NAND2_322 (.Y(N1318),.A(N715),.B(N1228));
INVX1 NOT1_323 (.Y(N1319),.A(N1158));
NAND2X1 NAND2_324 (.Y(N1322),.A(N628),.B(N1230));
NAND2X1 NAND2_325 (.Y(N1327),.A(N730),.B(N1238));
NAND2X1 NAND2_326 (.Y(N1328),.A(N733),.B(N1241));
INVX1 NOT1_327 (.Y(N1334),.A(N1162));
NAND2X1 NAND2_328 (.Y(N1344),.A(N1267),.B(N1160));
NAND2X1 NAND2_329 (.Y(N1345),.A(N1249),.B(N894));
INVX1 NOT1_330 (.Y(N1346),.A(N1249));
INVX1 NOT1_331 (.Y(N1348),.A(N1255));
INVX1 NOT1_332 (.Y(N1349),.A(N1252));
INVX1 NOT1_333 (.Y(N1350),.A(N1261));
INVX1 NOT1_334 (.Y(N1351),.A(N1258));
NAND2X1 NAND2_335 (.Y(N1352),.A(N1309),.B(N1206));
NAND2X1 NAND2_336 (.Y(N1355),.A(N1310),.B(N1208));
NAND2X1 NAND2_337 (.Y(N1358),.A(N1311),.B(N1210));
NAND2X1 NAND2_338 (.Y(N1361),.A(N1312),.B(N1212));
NAND2X1 NAND2_339 (.Y(N1364),.A(N1313),.B(N1214));
NAND2X1 NAND2_340 (.Y(N1367),.A(N1314),.B(N1216));
NAND2X1 NAND2_341 (.Y(N1370),.A(N1315),.B(N1221));
NAND2X1 NAND2_342 (.Y(N1373),.A(N1316),.B(N1224));
NAND2X1 NAND2_343 (.Y(N1376),.A(N1317),.B(N1226));
NAND2X1 NAND2_344 (.Y(N1379),.A(N1318),.B(N1229));
NAND2X1 NAND2_345 (.Y(N1383),.A(N1322),.B(N1231));
INVX1 NOT1_346 (.Y(N1386),.A(N1232));
NAND2X1 NAND2_347 (.Y(N1387),.A(N1232),.B(N990));
INVX1 NOT1_348 (.Y(N1388),.A(N1235));
NAND2X1 NAND2_349 (.Y(N1389),.A(N1235),.B(N993));
NAND2X1 NAND2_350 (.Y(N1390),.A(N1327),.B(N1239));
NAND2X1 NAND2_351 (.Y(N1393),.A(N1328),.B(N1242));
INVX1 NOT1_352 (.Y(N1396),.A(N1243));
NAND2X1 NAND2_353 (.Y(N1397),.A(N1243),.B(N1004));
INVX1 NOT1_354 (.Y(N1398),.A(N1246));
NAND2X1 NAND2_355 (.Y(N1399),.A(N1246),.B(N1007));
INVX1 NOT1_356 (.Y(N1409),.A(N1319));
NAND2X1 NAND2_357 (.Y(N1412),.A(N649),.B(N1346));
INVX1 NOT1_358 (.Y(N1413),.A(N1334));
BUFX1 BUFF1_359 (.Y(N1416),.A(N1264));
BUFX1 BUFF1_360 (.Y(N1419),.A(N1264));
NAND2X1 NAND2_361 (.Y(N1433),.A(N634),.B(N1386));
NAND2X1 NAND2_362 (.Y(N1434),.A(N637),.B(N1388));
NAND2X1 NAND2_363 (.Y(N1438),.A(N640),.B(N1396));
NAND2X1 NAND2_364 (.Y(N1439),.A(N646),.B(N1398));
INVX1 NOT1_365 (.Y(N1440),.A(N1344));
NAND2X1 NAND2_366 (.Y(N1443),.A(N1355),.B(N1148));
INVX1 NOT1_367 (.Y(N1444),.A(N1355));
NAND2X1 NAND2_368 (.Y(N1445),.A(N1352),.B(N1149));
INVX1 NOT1_369 (.Y(N1446),.A(N1352));
NAND2X1 NAND2_370 (.Y(N1447),.A(N1358),.B(N1151));
INVX1 NOT1_371 (.Y(N1448),.A(N1358));
NAND2X1 NAND2_372 (.Y(N1451),.A(N1361),.B(N1152));
INVX1 NOT1_373 (.Y(N1452),.A(N1361));
NAND2X1 NAND2_374 (.Y(N1453),.A(N1367),.B(N1153));
INVX1 NOT1_375 (.Y(N1454),.A(N1367));
NAND2X1 NAND2_376 (.Y(N1455),.A(N1364),.B(N1154));
INVX1 NOT1_377 (.Y(N1456),.A(N1364));
NAND2X1 NAND2_378 (.Y(N1457),.A(N1373),.B(N1156));
INVX1 NOT1_379 (.Y(N1458),.A(N1373));
NAND2X1 NAND2_380 (.Y(N1459),.A(N1379),.B(N1157));
INVX1 NOT1_381 (.Y(N1460),.A(N1379));
INVX1 NOT1_382 (.Y(N1461),.A(N1383));
NAND2X1 NAND2_383 (.Y(N1462),.A(N1393),.B(N1161));
INVX1 NOT1_384 (.Y(N1463),.A(N1393));
NAND2X1 NAND2_385 (.Y(N1464),.A(N1345),.B(N1412));
INVX1 NOT1_386 (.Y(N1468),.A(N1370));
NAND2X1 NAND2_387 (.Y(N1469),.A(N1370),.B(N1222));
INVX1 NOT1_388 (.Y(N1470),.A(N1376));
NAND2X1 NAND2_389 (.Y(N1471),.A(N1376),.B(N1227));
NAND2X1 NAND2_390 (.Y(N1472),.A(N1387),.B(N1433));
INVX1 NOT1_391 (.Y(N1475),.A(N1390));
NAND2X1 NAND2_392 (.Y(N1476),.A(N1390),.B(N1240));
NAND2X1 NAND2_393 (.Y(N1478),.A(N1389),.B(N1434));
NAND2X1 NAND2_394 (.Y(N1481),.A(N1399),.B(N1439));
NAND2X1 NAND2_395 (.Y(N1484),.A(N1397),.B(N1438));
NAND2X1 NAND2_396 (.Y(N1487),.A(N939),.B(N1444));
NAND2X1 NAND2_397 (.Y(N1488),.A(N935),.B(N1446));
NAND2X1 NAND2_398 (.Y(N1489),.A(N943),.B(N1448));
INVX1 NOT1_399 (.Y(N1490),.A(N1419));
INVX1 NOT1_400 (.Y(N1491),.A(N1416));
NAND2X1 NAND2_401 (.Y(N1492),.A(N947),.B(N1452));
NAND2X1 NAND2_402 (.Y(N1493),.A(N955),.B(N1454));
NAND2X1 NAND2_403 (.Y(N1494),.A(N951),.B(N1456));
NAND2X1 NAND2_404 (.Y(N1495),.A(N969),.B(N1458));
NAND2X1 NAND2_405 (.Y(N1496),.A(N977),.B(N1460));
NAND2X1 NAND2_406 (.Y(N1498),.A(N998),.B(N1463));
INVX1 NOT1_407 (.Y(N1499),.A(N1440));
NAND2X1 NAND2_408 (.Y(N1500),.A(N965),.B(N1468));
NAND2X1 NAND2_409 (.Y(N1501),.A(N973),.B(N1470));
NAND2X1 NAND2_410 (.Y(N1504),.A(N994),.B(N1475));
INVX1 NOT1_411 (.Y(N1510),.A(N1464));
NAND2X1 NAND2_412 (.Y(N1513),.A(N1443),.B(N1487));
NAND2X1 NAND2_413 (.Y(N1514),.A(N1445),.B(N1488));
NAND2X1 NAND2_414 (.Y(N1517),.A(N1447),.B(N1489));
NAND2X1 NAND2_415 (.Y(N1520),.A(N1451),.B(N1492));
NAND2X1 NAND2_416 (.Y(N1521),.A(N1453),.B(N1493));
NAND2X1 NAND2_417 (.Y(N1522),.A(N1455),.B(N1494));
NAND2X1 NAND2_418 (.Y(N1526),.A(N1457),.B(N1495));
NAND2X1 NAND2_419 (.Y(N1527),.A(N1459),.B(N1496));
INVX1 NOT1_420 (.Y(N1528),.A(N1472));
NAND2X1 NAND2_421 (.Y(N1529),.A(N1462),.B(N1498));
INVX1 NOT1_422 (.Y(N1530),.A(N1478));
INVX1 NOT1_423 (.Y(N1531),.A(N1481));
INVX1 NOT1_424 (.Y(N1532),.A(N1484));
NAND2X1 NAND2_425 (.Y(N1534),.A(N1471),.B(N1501));
NAND2X1 NAND2_426 (.Y(N1537),.A(N1469),.B(N1500));
NAND2X1 NAND2_427 (.Y(N1540),.A(N1476),.B(N1504));
INVX1 NOT1_428 (.Y(N1546),.A(N1513));
INVX1 NOT1_429 (.Y(N1554),.A(N1521));
INVX1 NOT1_430 (.Y(N1557),.A(N1526));
INVX1 NOT1_431 (.Y(N1561),.A(N1520));
NAND2X1 NAND2_432 (.Y(N1567),.A(N1484),.B(N1531));
NAND2X1 NAND2_433 (.Y(N1568),.A(N1481),.B(N1532));
INVX1 NOT1_434 (.Y(N1569),.A(N1510));
INVX1 NOT1_435 (.Y(N1571),.A(N1527));
INVX1 NOT1_436 (.Y(N1576),.A(N1529));
BUFX1 BUFF1_437 (.Y(N1588),.A(N1522));
INVX1 NOT1_438 (.Y(N1591),.A(N1534));
INVX1 NOT1_439 (.Y(N1593),.A(N1537));
NAND2X1 NAND2_440 (.Y(N1594),.A(N1540),.B(N1530));
INVX1 NOT1_441 (.Y(N1595),.A(N1540));
NAND2X1 NAND2_442 (.Y(N1596),.A(N1567),.B(N1568));
BUFX1 BUFF1_443 (.Y(N1600),.A(N1517));
BUFX1 BUFF1_444 (.Y(N1603),.A(N1517));
BUFX1 BUFF1_445 (.Y(N1606),.A(N1522));
BUFX1 BUFF1_446 (.Y(N1609),.A(N1522));
BUFX1 BUFF1_447 (.Y(N1612),.A(N1514));
BUFX1 BUFF1_448 (.Y(N1615),.A(N1514));
BUFX1 BUFF1_449 (.Y(N1620),.A(N1557));
BUFX1 BUFF1_450 (.Y(N1623),.A(N1554));
INVX1 NOT1_451 (.Y(N1635),.A(N1571));
NAND2X1 NAND2_452 (.Y(N1636),.A(N1478),.B(N1595));
NAND2X1 NAND2_453 (.Y(N1638),.A(N1576),.B(N1569));
INVX1 NOT1_454 (.Y(N1639),.A(N1576));
BUFX1 BUFF1_455 (.Y(N1640),.A(N1561));
BUFX1 BUFF1_456 (.Y(N1643),.A(N1561));
BUFX1 BUFF1_457 (.Y(N1647),.A(N1546));
BUFX1 BUFF1_458 (.Y(N1651),.A(N1546));
BUFX1 BUFF1_459 (.Y(N1658),.A(N1554));
BUFX1 BUFF1_460 (.Y(N1661),.A(N1557));
BUFX1 BUFF1_461 (.Y(N1664),.A(N1557));
NAND2X1 NAND2_462 (.Y(N1671),.A(N1596),.B(N893));
INVX1 NOT1_463 (.Y(N1672),.A(N1596));
INVX1 NOT1_464 (.Y(N1675),.A(N1600));
INVX1 NOT1_465 (.Y(N1677),.A(N1603));
NAND2X1 NAND2_466 (.Y(N1678),.A(N1606),.B(N1217));
INVX1 NOT1_467 (.Y(N1679),.A(N1606));
NAND2X1 NAND2_468 (.Y(N1680),.A(N1609),.B(N1219));
INVX1 NOT1_469 (.Y(N1681),.A(N1609));
INVX1 NOT1_470 (.Y(N1682),.A(N1612));
INVX1 NOT1_471 (.Y(N1683),.A(N1615));
NAND2X1 NAND2_472 (.Y(N1685),.A(N1594),.B(N1636));
NAND2X1 NAND2_473 (.Y(N1688),.A(N1510),.B(N1639));
BUFX1 BUFF1_474 (.Y(N1697),.A(N1588));
BUFX1 BUFF1_475 (.Y(N1701),.A(N1588));
NAND2X1 NAND2_476 (.Y(N1706),.A(N643),.B(N1672));
INVX1 NOT1_477 (.Y(N1707),.A(N1643));
NAND2X1 NAND2_478 (.Y(N1708),.A(N1647),.B(N1675));
INVX1 NOT1_479 (.Y(N1709),.A(N1647));
NAND2X1 NAND2_480 (.Y(N1710),.A(N1651),.B(N1677));
INVX1 NOT1_481 (.Y(N1711),.A(N1651));
NAND2X1 NAND2_482 (.Y(N1712),.A(N1028),.B(N1679));
NAND2X1 NAND2_483 (.Y(N1713),.A(N1031),.B(N1681));
BUFX1 BUFF1_484 (.Y(N1714),.A(N1620));
BUFX1 BUFF1_485 (.Y(N1717),.A(N1620));
NAND2X1 NAND2_486 (.Y(N1720),.A(N1658),.B(N1593));
INVX1 NOT1_487 (.Y(N1721),.A(N1658));
NAND2X1 NAND2_488 (.Y(N1723),.A(N1638),.B(N1688));
INVX1 NOT1_489 (.Y(N1727),.A(N1661));
INVX1 NOT1_490 (.Y(N1728),.A(N1640));
INVX1 NOT1_491 (.Y(N1730),.A(N1664));
BUFX1 BUFF1_492 (.Y(N1731),.A(N1623));
BUFX1 BUFF1_493 (.Y(N1734),.A(N1623));
NAND2X1 NAND2_494 (.Y(N1740),.A(N1685),.B(N1528));
INVX1 NOT1_495 (.Y(N1741),.A(N1685));
NAND2X1 NAND2_496 (.Y(N1742),.A(N1671),.B(N1706));
NAND2X1 NAND2_497 (.Y(N1746),.A(N1600),.B(N1709));
NAND2X1 NAND2_498 (.Y(N1747),.A(N1603),.B(N1711));
NAND2X1 NAND2_499 (.Y(N1748),.A(N1678),.B(N1712));
NAND2X1 NAND2_500 (.Y(N1751),.A(N1680),.B(N1713));
NAND2X1 NAND2_501 (.Y(N1759),.A(N1537),.B(N1721));
INVX1 NOT1_502 (.Y(N1761),.A(N1697));
NAND2X1 NAND2_503 (.Y(N1762),.A(N1697),.B(N1727));
INVX1 NOT1_504 (.Y(N1763),.A(N1701));
NAND2X1 NAND2_505 (.Y(N1764),.A(N1701),.B(N1730));
INVX1 NOT1_506 (.Y(N1768),.A(N1717));
NAND2X1 NAND2_507 (.Y(N1769),.A(N1472),.B(N1741));
NAND2X1 NAND2_508 (.Y(N1772),.A(N1723),.B(N1413));
INVX1 NOT1_509 (.Y(N1773),.A(N1723));
NAND2X1 NAND2_510 (.Y(N1774),.A(N1708),.B(N1746));
NAND2X1 NAND2_511 (.Y(N1777),.A(N1710),.B(N1747));
INVX1 NOT1_512 (.Y(N1783),.A(N1731));
NAND2X1 NAND2_513 (.Y(N1784),.A(N1731),.B(N1682));
INVX1 NOT1_514 (.Y(N1785),.A(N1714));
INVX1 NOT1_515 (.Y(N1786),.A(N1734));
NAND2X1 NAND2_516 (.Y(N1787),.A(N1734),.B(N1683));
NAND2X1 NAND2_517 (.Y(N1788),.A(N1720),.B(N1759));
NAND2X1 NAND2_518 (.Y(N1791),.A(N1661),.B(N1761));
NAND2X1 NAND2_519 (.Y(N1792),.A(N1664),.B(N1763));
NAND2X1 NAND2_520 (.Y(N1795),.A(N1751),.B(N1155));
INVX1 NOT1_521 (.Y(N1796),.A(N1751));
NAND2X1 NAND2_522 (.Y(N1798),.A(N1740),.B(N1769));
NAND2X1 NAND2_523 (.Y(N1801),.A(N1334),.B(N1773));
NAND2X1 NAND2_524 (.Y(N1802),.A(N1742),.B(N290));
INVX1 NOT1_525 (.Y(N1807),.A(N1748));
NAND2X1 NAND2_526 (.Y(N1808),.A(N1748),.B(N1218));
NAND2X1 NAND2_527 (.Y(N1809),.A(N1612),.B(N1783));
NAND2X1 NAND2_528 (.Y(N1810),.A(N1615),.B(N1786));
NAND2X1 NAND2_529 (.Y(N1812),.A(N1791),.B(N1762));
NAND2X1 NAND2_530 (.Y(N1815),.A(N1792),.B(N1764));
BUFX1 BUFF1_531 (.Y(N1818),.A(N1742));
NAND2X1 NAND2_532 (.Y(N1821),.A(N1777),.B(N1490));
INVX1 NOT1_533 (.Y(N1822),.A(N1777));
NAND2X1 NAND2_534 (.Y(N1823),.A(N1774),.B(N1491));
INVX1 NOT1_535 (.Y(N1824),.A(N1774));
NAND2X1 NAND2_536 (.Y(N1825),.A(N962),.B(N1796));
NAND2X1 NAND2_537 (.Y(N1826),.A(N1788),.B(N1409));
INVX1 NOT1_538 (.Y(N1827),.A(N1788));
NAND2X1 NAND2_539 (.Y(N1830),.A(N1772),.B(N1801));
NAND2X1 NAND2_540 (.Y(N1837),.A(N959),.B(N1807));
NAND2X1 NAND2_541 (.Y(N1838),.A(N1809),.B(N1784));
NAND2X1 NAND2_542 (.Y(N1841),.A(N1810),.B(N1787));
NAND2X1 NAND2_543 (.Y(N1848),.A(N1419),.B(N1822));
NAND2X1 NAND2_544 (.Y(N1849),.A(N1416),.B(N1824));
NAND2X1 NAND2_545 (.Y(N1850),.A(N1795),.B(N1825));
NAND2X1 NAND2_546 (.Y(N1852),.A(N1319),.B(N1827));
NAND2X1 NAND2_547 (.Y(N1855),.A(N1815),.B(N1707));
INVX1 NOT1_548 (.Y(N1856),.A(N1815));
INVX1 NOT1_549 (.Y(N1857),.A(N1818));
NAND2X1 NAND2_550 (.Y(N1858),.A(N1798),.B(N290));
INVX1 NOT1_551 (.Y(N1864),.A(N1812));
NAND2X1 NAND2_552 (.Y(N1865),.A(N1812),.B(N1728));
BUFX1 BUFF1_553 (.Y(N1866),.A(N1798));
BUFX1 BUFF1_554 (.Y(N1869),.A(N1802));
BUFX1 BUFF1_555 (.Y(N1872),.A(N1802));
NAND2X1 NAND2_556 (.Y(N1875),.A(N1808),.B(N1837));
NAND2X1 NAND2_557 (.Y(N1878),.A(N1821),.B(N1848));
NAND2X1 NAND2_558 (.Y(N1879),.A(N1823),.B(N1849));
NAND2X1 NAND2_559 (.Y(N1882),.A(N1841),.B(N1768));
INVX1 NOT1_560 (.Y(N1883),.A(N1841));
NAND2X1 NAND2_561 (.Y(N1884),.A(N1826),.B(N1852));
NAND2X1 NAND2_562 (.Y(N1885),.A(N1643),.B(N1856));
NAND2X1 NAND2_563 (.Y(N1889),.A(N1830),.B(N290));
INVX1 NOT1_564 (.Y(N1895),.A(N1838));
NAND2X1 NAND2_565 (.Y(N1896),.A(N1838),.B(N1785));
NAND2X1 NAND2_566 (.Y(N1897),.A(N1640),.B(N1864));
INVX1 NOT1_567 (.Y(N1898),.A(N1850));
BUFX1 BUFF1_568 (.Y(N1902),.A(N1830));
INVX1 NOT1_569 (.Y(N1910),.A(N1878));
NAND2X1 NAND2_570 (.Y(N1911),.A(N1717),.B(N1883));
INVX1 NOT1_571 (.Y(N1912),.A(N1884));
NAND2X1 NAND2_572 (.Y(N1913),.A(N1855),.B(N1885));
INVX1 NOT1_573 (.Y(N1915),.A(N1866));
NAND2X1 NAND2_574 (.Y(N1919),.A(N1872),.B(N919));
INVX1 NOT1_575 (.Y(N1920),.A(N1872));
NAND2X1 NAND2_576 (.Y(N1921),.A(N1869),.B(N920));
INVX1 NOT1_577 (.Y(N1922),.A(N1869));
INVX1 NOT1_578 (.Y(N1923),.A(N1875));
NAND2X1 NAND2_579 (.Y(N1924),.A(N1714),.B(N1895));
BUFX1 BUFF1_580 (.Y(N1927),.A(N1858));
BUFX1 BUFF1_581 (.Y(N1930),.A(N1858));
NAND2X1 NAND2_582 (.Y(N1933),.A(N1865),.B(N1897));
NAND2X1 NAND2_583 (.Y(N1936),.A(N1882),.B(N1911));
INVX1 NOT1_584 (.Y(N1937),.A(N1898));
INVX1 NOT1_585 (.Y(N1938),.A(N1902));
NAND2X1 NAND2_586 (.Y(N1941),.A(N679),.B(N1920));
NAND2X1 NAND2_587 (.Y(N1942),.A(N676),.B(N1922));
BUFX1 BUFF1_588 (.Y(N1944),.A(N1879));
INVX1 NOT1_589 (.Y(N1947),.A(N1913));
BUFX1 BUFF1_590 (.Y(N1950),.A(N1889));
BUFX1 BUFF1_591 (.Y(N1953),.A(N1889));
BUFX1 BUFF1_592 (.Y(N1958),.A(N1879));
NAND2X1 NAND2_593 (.Y(N1961),.A(N1896),.B(N1924));
AND2X1 AND2_594 (.Y(N1965),.A(N1910),.B(N601));
AND2X1 AND2_595 (.Y(N1968),.A(N602),.B(N1912));
NAND2X1 NAND2_596 (.Y(N1975),.A(N1930),.B(N917));
INVX1 NOT1_597 (.Y(N1976),.A(N1930));
NAND2X1 NAND2_598 (.Y(N1977),.A(N1927),.B(N918));
INVX1 NOT1_599 (.Y(N1978),.A(N1927));
NAND2X1 NAND2_600 (.Y(N1979),.A(N1919),.B(N1941));
NAND2X1 NAND2_601 (.Y(N1980),.A(N1921),.B(N1942));
INVX1 NOT1_602 (.Y(N1985),.A(N1933));
INVX1 NOT1_603 (.Y(N1987),.A(N1936));
INVX1 NOT1_604 (.Y(N1999),.A(N1944));
NAND2X1 NAND2_605 (.Y(N2000),.A(N1944),.B(N1937));
INVX1 NOT1_606 (.Y(N2002),.A(N1947));
NAND2X1 NAND2_607 (.Y(N2003),.A(N1947),.B(N1499));
NAND2X1 NAND2_608 (.Y(N2004),.A(N1953),.B(N1350));
INVX1 NOT1_609 (.Y(N2005),.A(N1953));
NAND2X1 NAND2_610 (.Y(N2006),.A(N1950),.B(N1351));
INVX1 NOT1_611 (.Y(N2007),.A(N1950));
NAND2X1 NAND2_612 (.Y(N2008),.A(N673),.B(N1976));
NAND2X1 NAND2_613 (.Y(N2009),.A(N670),.B(N1978));
INVX1 NOT1_614 (.Y(N2012),.A(N1979));
INVX1 NOT1_615 (.Y(N2013),.A(N1958));
NAND2X1 NAND2_616 (.Y(N2014),.A(N1958),.B(N1923));
INVX1 NOT1_617 (.Y(N2015),.A(N1961));
NAND2X1 NAND2_618 (.Y(N2016),.A(N1961),.B(N1635));
INVX1 NOT1_619 (.Y(N2018),.A(N1965));
INVX1 NOT1_620 (.Y(N2019),.A(N1968));
NAND2X1 NAND2_621 (.Y(N2020),.A(N1898),.B(N1999));
INVX1 NOT1_622 (.Y(N2021),.A(N1987));
NAND2X1 NAND2_623 (.Y(N2022),.A(N1987),.B(N1591));
NAND2X1 NAND2_624 (.Y(N2023),.A(N1440),.B(N2002));
NAND2X1 NAND2_625 (.Y(N2024),.A(N1261),.B(N2005));
NAND2X1 NAND2_626 (.Y(N2025),.A(N1258),.B(N2007));
NAND2X1 NAND2_627 (.Y(N2026),.A(N1975),.B(N2008));
NAND2X1 NAND2_628 (.Y(N2027),.A(N1977),.B(N2009));
INVX1 NOT1_629 (.Y(N2030),.A(N1980));
BUFX1 BUFF1_630 (.Y(N2033),.A(N1980));
NAND2X1 NAND2_631 (.Y(N2036),.A(N1875),.B(N2013));
NAND2X1 NAND2_632 (.Y(N2037),.A(N1571),.B(N2015));
NAND2X1 NAND2_633 (.Y(N2038),.A(N2020),.B(N2000));
NAND2X1 NAND2_634 (.Y(N2039),.A(N1534),.B(N2021));
NAND2X1 NAND2_635 (.Y(N2040),.A(N2023),.B(N2003));
NAND2X1 NAND2_636 (.Y(N2041),.A(N2004),.B(N2024));
NAND2X1 NAND2_637 (.Y(N2042),.A(N2006),.B(N2025));
INVX1 NOT1_638 (.Y(N2047),.A(N2026));
NAND2X1 NAND2_639 (.Y(N2052),.A(N2036),.B(N2014));
NAND2X1 NAND2_640 (.Y(N2055),.A(N2037),.B(N2016));
INVX1 NOT1_641 (.Y(N2060),.A(N2038));
NAND2X1 NAND2_642 (.Y(N2061),.A(N2039),.B(N2022));
NAND2X1 NAND2_643 (.Y(N2062),.A(N2040),.B(N290));
INVX1 NOT1_644 (.Y(N2067),.A(N2041));
INVX1 NOT1_645 (.Y(N2068),.A(N2027));
BUFX1 BUFF1_646 (.Y(N2071),.A(N2027));
INVX1 NOT1_647 (.Y(N2076),.A(N2052));
INVX1 NOT1_648 (.Y(N2077),.A(N2055));
NAND2X1 NAND2_649 (.Y(N2078),.A(N2060),.B(N290));
NAND2X1 NAND2_650 (.Y(N2081),.A(N2061),.B(N290));
INVX1 NOT1_651 (.Y(N2086),.A(N2042));
BUFX1 BUFF1_652 (.Y(N2089),.A(N2042));
AND2X1 AND2_653 (.Y(N2104),.A(N2030),.B(N2068));
AND2X1 AND2_654 (.Y(N2119),.A(N2033),.B(N2068));
AND2X1 AND2_655 (.Y(N2129),.A(N2030),.B(N2071));
AND2X1 AND2_656 (.Y(N2143),.A(N2033),.B(N2071));
BUFX1 BUFF1_657 (.Y(N2148),.A(N2062));
BUFX1 BUFF1_658 (.Y(N2151),.A(N2062));
BUFX1 BUFF1_659 (.Y(N2196),.A(N2078));
BUFX1 BUFF1_660 (.Y(N2199),.A(N2078));
BUFX1 BUFF1_661 (.Y(N2202),.A(N2081));
BUFX1 BUFF1_662 (.Y(N2205),.A(N2081));
NAND2X1 NAND2_663 (.Y(N2214),.A(N2151),.B(N915));
INVX1 NOT1_664 (.Y(N2215),.A(N2151));
NAND2X1 NAND2_665 (.Y(N2216),.A(N2148),.B(N916));
INVX1 NOT1_666 (.Y(N2217),.A(N2148));
NAND2X1 NAND2_667 (.Y(N2222),.A(N2199),.B(N1348));
INVX1 NOT1_668 (.Y(N2223),.A(N2199));
NAND2X1 NAND2_669 (.Y(N2224),.A(N2196),.B(N1349));
INVX1 NOT1_670 (.Y(N2225),.A(N2196));
NAND2X1 NAND2_671 (.Y(N2226),.A(N2205),.B(N913));
INVX1 NOT1_672 (.Y(N2227),.A(N2205));
NAND2X1 NAND2_673 (.Y(N2228),.A(N2202),.B(N914));
INVX1 NOT1_674 (.Y(N2229),.A(N2202));
NAND2X1 NAND2_675 (.Y(N2230),.A(N667),.B(N2215));
NAND2X1 NAND2_676 (.Y(N2231),.A(N664),.B(N2217));
NAND2X1 NAND2_677 (.Y(N2232),.A(N1255),.B(N2223));
NAND2X1 NAND2_678 (.Y(N2233),.A(N1252),.B(N2225));
NAND2X1 NAND2_679 (.Y(N2234),.A(N661),.B(N2227));
NAND2X1 NAND2_680 (.Y(N2235),.A(N658),.B(N2229));
NAND2X1 NAND2_681 (.Y(N2236),.A(N2214),.B(N2230));
NAND2X1 NAND2_682 (.Y(N2237),.A(N2216),.B(N2231));
NAND2X1 NAND2_683 (.Y(N2240),.A(N2222),.B(N2232));
NAND2X1 NAND2_684 (.Y(N2241),.A(N2224),.B(N2233));
NAND2X1 NAND2_685 (.Y(N2244),.A(N2226),.B(N2234));
NAND2X1 NAND2_686 (.Y(N2245),.A(N2228),.B(N2235));
INVX1 NOT1_687 (.Y(N2250),.A(N2236));
INVX1 NOT1_688 (.Y(N2253),.A(N2240));
INVX1 NOT1_689 (.Y(N2256),.A(N2244));
INVX1 NOT1_690 (.Y(N2257),.A(N2237));
BUFX1 BUFF1_691 (.Y(N2260),.A(N2237));
INVX1 NOT1_692 (.Y(N2263),.A(N2241));
AND2X1 AND2_693 (.Y(N2266),.A(N1164),.B(N2241));
INVX1 NOT1_694 (.Y(N2269),.A(N2245));
AND2X1 AND2_695 (.Y(N2272),.A(N1168),.B(N2245));
AND2X1 AND_tmp19 (.Y(ttmp19),.A(N2253),.B(N903));
AND2X1 AND_tmp20 (.Y(ttmp20),.A(N2067),.B(ttmp19));
AND2X1 AND_tmp21 (.Y(ttmp21),.A(N2012),.B(ttmp20));
AND2X1 AND_tmp22 (.Y(ttmp22),.A(N2047),.B(ttmp21));
AND2X1 AND_tmp23 (.Y(ttmp23),.A(N2250),.B(ttmp22));
AND2X1 AND_tmp24 (.Y(ttmp24),.A(N899),.B(ttmp23));
NAND2X1 NAND_tmp25 (.Y(N2279),.A(N2256),.B(ttmp24));
BUFX1 BUFF1_697 (.Y(N2286),.A(N2266));
BUFX1 BUFF1_698 (.Y(N2297),.A(N2266));
BUFX1 BUFF1_699 (.Y(N2315),.A(N2272));
BUFX1 BUFF1_700 (.Y(N2326),.A(N2272));
AND2X1 AND2_701 (.Y(N2340),.A(N2086),.B(N2257));
AND2X1 AND2_702 (.Y(N2353),.A(N2089),.B(N2257));
AND2X1 AND2_703 (.Y(N2361),.A(N2086),.B(N2260));
AND2X1 AND2_704 (.Y(N2375),.A(N2089),.B(N2260));
AND2X1 AND_tmp26 (.Y(ttmp26),.A(N313),.B(N313));
AND2X1 AND_tmp27 (.Y(ttmp27),.A(N338),.B(ttmp26));
AND2X1 AND_tmp28 (.Y(N2384),.A(N2279),.B(ttmp27));
AND2X1 AND2_706 (.Y(N2385),.A(N1163),.B(N2263));
AND2X1 AND2_707 (.Y(N2386),.A(N1164),.B(N2263));
AND2X1 AND2_708 (.Y(N2426),.A(N1167),.B(N2269));
AND2X1 AND2_709 (.Y(N2427),.A(N1168),.B(N2269));
AND2X1 AND_tmp29 (.Y(ttmp29),.A(N2104),.B(N1171));
AND2X1 AND_tmp30 (.Y(ttmp30),.A(N2286),.B(ttmp29));
AND2X1 AND_tmp31 (.Y(ttmp31),.A(N2315),.B(ttmp30));
NAND2X1 NAND_tmp32 (.Y(N2537),.A(N2361),.B(ttmp31));
AND2X1 AND_tmp33 (.Y(ttmp33),.A(N2129),.B(N1171));
AND2X1 AND_tmp34 (.Y(ttmp34),.A(N2286),.B(ttmp33));
AND2X1 AND_tmp35 (.Y(ttmp35),.A(N2315),.B(ttmp34));
NAND2X1 NAND_tmp36 (.Y(N2540),.A(N2340),.B(ttmp35));
AND2X1 AND_tmp37 (.Y(ttmp37),.A(N2119),.B(N1171));
AND2X1 AND_tmp38 (.Y(ttmp38),.A(N2286),.B(ttmp37));
AND2X1 AND_tmp39 (.Y(ttmp39),.A(N2315),.B(ttmp38));
NAND2X1 NAND_tmp40 (.Y(N2543),.A(N2340),.B(ttmp39));
AND2X1 AND_tmp41 (.Y(ttmp41),.A(N2104),.B(N1171));
AND2X1 AND_tmp42 (.Y(ttmp42),.A(N2286),.B(ttmp41));
AND2X1 AND_tmp43 (.Y(ttmp43),.A(N2315),.B(ttmp42));
NAND2X1 NAND_tmp44 (.Y(N2546),.A(N2353),.B(ttmp43));
AND2X1 AND_tmp45 (.Y(ttmp45),.A(N2119),.B(N1188));
AND2X1 AND_tmp46 (.Y(ttmp46),.A(N2297),.B(ttmp45));
AND2X1 AND_tmp47 (.Y(ttmp47),.A(N2315),.B(ttmp46));
NAND2X1 NAND_tmp48 (.Y(N2549),.A(N2375),.B(ttmp47));
AND2X1 AND_tmp49 (.Y(ttmp49),.A(N2143),.B(N1188));
AND2X1 AND_tmp50 (.Y(ttmp50),.A(N2297),.B(ttmp49));
AND2X1 AND_tmp51 (.Y(ttmp51),.A(N2326),.B(ttmp50));
NAND2X1 NAND_tmp52 (.Y(N2552),.A(N2361),.B(ttmp51));
AND2X1 AND_tmp53 (.Y(ttmp53),.A(N2129),.B(N1188));
AND2X1 AND_tmp54 (.Y(ttmp54),.A(N2297),.B(ttmp53));
AND2X1 AND_tmp55 (.Y(ttmp55),.A(N2326),.B(ttmp54));
NAND2X1 NAND_tmp56 (.Y(N2555),.A(N2375),.B(ttmp55));
AND2X1 AND_tmp57 (.Y(ttmp57),.A(N2104),.B(N1171));
AND2X1 AND_tmp58 (.Y(ttmp58),.A(N2286),.B(ttmp57));
AND2X1 AND_tmp59 (.Y(ttmp59),.A(N2315),.B(ttmp58));
AND2X1 AND_tmp60 (.Y(N2558),.A(N2361),.B(ttmp59));
AND2X1 AND_tmp61 (.Y(ttmp61),.A(N2129),.B(N1171));
AND2X1 AND_tmp62 (.Y(ttmp62),.A(N2286),.B(ttmp61));
AND2X1 AND_tmp63 (.Y(ttmp63),.A(N2315),.B(ttmp62));
AND2X1 AND_tmp64 (.Y(N2561),.A(N2340),.B(ttmp63));
AND2X1 AND_tmp65 (.Y(ttmp65),.A(N2119),.B(N1171));
AND2X1 AND_tmp66 (.Y(ttmp66),.A(N2286),.B(ttmp65));
AND2X1 AND_tmp67 (.Y(ttmp67),.A(N2315),.B(ttmp66));
AND2X1 AND_tmp68 (.Y(N2564),.A(N2340),.B(ttmp67));
AND2X1 AND_tmp69 (.Y(ttmp69),.A(N2104),.B(N1171));
AND2X1 AND_tmp70 (.Y(ttmp70),.A(N2286),.B(ttmp69));
AND2X1 AND_tmp71 (.Y(ttmp71),.A(N2315),.B(ttmp70));
AND2X1 AND_tmp72 (.Y(N2567),.A(N2353),.B(ttmp71));
AND2X1 AND_tmp73 (.Y(ttmp73),.A(N2119),.B(N1188));
AND2X1 AND_tmp74 (.Y(ttmp74),.A(N2297),.B(ttmp73));
AND2X1 AND_tmp75 (.Y(ttmp75),.A(N2315),.B(ttmp74));
AND2X1 AND_tmp76 (.Y(N2570),.A(N2375),.B(ttmp75));
AND2X1 AND_tmp77 (.Y(ttmp77),.A(N2143),.B(N1188));
AND2X1 AND_tmp78 (.Y(ttmp78),.A(N2297),.B(ttmp77));
AND2X1 AND_tmp79 (.Y(ttmp79),.A(N2326),.B(ttmp78));
AND2X1 AND_tmp80 (.Y(N2573),.A(N2361),.B(ttmp79));
AND2X1 AND_tmp81 (.Y(ttmp81),.A(N2129),.B(N1188));
AND2X1 AND_tmp82 (.Y(ttmp82),.A(N2297),.B(ttmp81));
AND2X1 AND_tmp83 (.Y(ttmp83),.A(N2326),.B(ttmp82));
AND2X1 AND_tmp84 (.Y(N2576),.A(N2375),.B(ttmp83));
AND2X1 AND_tmp85 (.Y(ttmp85),.A(N2129),.B(N1171));
AND2X1 AND_tmp86 (.Y(ttmp86),.A(N2286),.B(ttmp85));
AND2X1 AND_tmp87 (.Y(ttmp87),.A(N2427),.B(ttmp86));
NAND2X1 NAND_tmp88 (.Y(N2594),.A(N2361),.B(ttmp87));
AND2X1 AND_tmp89 (.Y(ttmp89),.A(N2119),.B(N1171));
AND2X1 AND_tmp90 (.Y(ttmp90),.A(N2297),.B(ttmp89));
AND2X1 AND_tmp91 (.Y(ttmp91),.A(N2427),.B(ttmp90));
NAND2X1 NAND_tmp92 (.Y(N2597),.A(N2361),.B(ttmp91));
AND2X1 AND_tmp93 (.Y(ttmp93),.A(N2104),.B(N1171));
AND2X1 AND_tmp94 (.Y(ttmp94),.A(N2297),.B(ttmp93));
AND2X1 AND_tmp95 (.Y(ttmp95),.A(N2427),.B(ttmp94));
NAND2X1 NAND_tmp96 (.Y(N2600),.A(N2375),.B(ttmp95));
AND2X1 AND_tmp97 (.Y(ttmp97),.A(N2143),.B(N1171));
AND2X1 AND_tmp98 (.Y(ttmp98),.A(N2297),.B(ttmp97));
AND2X1 AND_tmp99 (.Y(ttmp99),.A(N2427),.B(ttmp98));
NAND2X1 NAND_tmp100 (.Y(N2603),.A(N2340),.B(ttmp99));
AND2X1 AND_tmp101 (.Y(ttmp101),.A(N2129),.B(N1188));
AND2X1 AND_tmp102 (.Y(ttmp102),.A(N2297),.B(ttmp101));
AND2X1 AND_tmp103 (.Y(ttmp103),.A(N2427),.B(ttmp102));
NAND2X1 NAND_tmp104 (.Y(N2606),.A(N2353),.B(ttmp103));
AND2X1 AND_tmp105 (.Y(ttmp105),.A(N2129),.B(N1188));
AND2X1 AND_tmp106 (.Y(ttmp106),.A(N2386),.B(ttmp105));
AND2X1 AND_tmp107 (.Y(ttmp107),.A(N2326),.B(ttmp106));
NAND2X1 NAND_tmp108 (.Y(N2611),.A(N2361),.B(ttmp107));
AND2X1 AND_tmp109 (.Y(ttmp109),.A(N2119),.B(N1188));
AND2X1 AND_tmp110 (.Y(ttmp110),.A(N2386),.B(ttmp109));
AND2X1 AND_tmp111 (.Y(ttmp111),.A(N2326),.B(ttmp110));
NAND2X1 NAND_tmp112 (.Y(N2614),.A(N2361),.B(ttmp111));
AND2X1 AND_tmp113 (.Y(ttmp113),.A(N2104),.B(N1188));
AND2X1 AND_tmp114 (.Y(ttmp114),.A(N2386),.B(ttmp113));
AND2X1 AND_tmp115 (.Y(ttmp115),.A(N2326),.B(ttmp114));
NAND2X1 NAND_tmp116 (.Y(N2617),.A(N2375),.B(ttmp115));
AND2X1 AND_tmp117 (.Y(ttmp117),.A(N2129),.B(N1188));
AND2X1 AND_tmp118 (.Y(ttmp118),.A(N2386),.B(ttmp117));
AND2X1 AND_tmp119 (.Y(ttmp119),.A(N2326),.B(ttmp118));
NAND2X1 NAND_tmp120 (.Y(N2620),.A(N2353),.B(ttmp119));
AND2X1 AND_tmp121 (.Y(ttmp121),.A(N2104),.B(N926));
AND2X1 AND_tmp122 (.Y(ttmp122),.A(N2297),.B(ttmp121));
AND2X1 AND_tmp123 (.Y(ttmp123),.A(N2427),.B(ttmp122));
NAND2X1 NAND_tmp124 (.Y(N2627),.A(N2340),.B(ttmp123));
AND2X1 AND_tmp125 (.Y(ttmp125),.A(N2104),.B(N926));
AND2X1 AND_tmp126 (.Y(ttmp126),.A(N2386),.B(ttmp125));
AND2X1 AND_tmp127 (.Y(ttmp127),.A(N2326),.B(ttmp126));
NAND2X1 NAND_tmp128 (.Y(N2628),.A(N2340),.B(ttmp127));
AND2X1 AND_tmp129 (.Y(ttmp129),.A(N2104),.B(N926));
AND2X1 AND_tmp130 (.Y(ttmp130),.A(N2386),.B(ttmp129));
AND2X1 AND_tmp131 (.Y(ttmp131),.A(N2427),.B(ttmp130));
NAND2X1 NAND_tmp132 (.Y(N2629),.A(N2361),.B(ttmp131));
AND2X1 AND_tmp133 (.Y(ttmp133),.A(N2129),.B(N926));
AND2X1 AND_tmp134 (.Y(ttmp134),.A(N2386),.B(ttmp133));
AND2X1 AND_tmp135 (.Y(ttmp135),.A(N2427),.B(ttmp134));
NAND2X1 NAND_tmp136 (.Y(N2630),.A(N2340),.B(ttmp135));
AND2X1 AND_tmp137 (.Y(ttmp137),.A(N2119),.B(N926));
AND2X1 AND_tmp138 (.Y(ttmp138),.A(N2386),.B(ttmp137));
AND2X1 AND_tmp139 (.Y(ttmp139),.A(N2427),.B(ttmp138));
NAND2X1 NAND_tmp140 (.Y(N2631),.A(N2340),.B(ttmp139));
AND2X1 AND_tmp141 (.Y(ttmp141),.A(N2104),.B(N926));
AND2X1 AND_tmp142 (.Y(ttmp142),.A(N2386),.B(ttmp141));
AND2X1 AND_tmp143 (.Y(ttmp143),.A(N2427),.B(ttmp142));
NAND2X1 NAND_tmp144 (.Y(N2632),.A(N2353),.B(ttmp143));
AND2X1 AND_tmp145 (.Y(ttmp145),.A(N2104),.B(N926));
AND2X1 AND_tmp146 (.Y(ttmp146),.A(N2386),.B(ttmp145));
AND2X1 AND_tmp147 (.Y(ttmp147),.A(N2426),.B(ttmp146));
NAND2X1 NAND_tmp148 (.Y(N2633),.A(N2340),.B(ttmp147));
AND2X1 AND_tmp149 (.Y(ttmp149),.A(N2104),.B(N926));
AND2X1 AND_tmp150 (.Y(ttmp150),.A(N2385),.B(ttmp149));
AND2X1 AND_tmp151 (.Y(ttmp151),.A(N2427),.B(ttmp150));
NAND2X1 NAND_tmp152 (.Y(N2634),.A(N2340),.B(ttmp151));
AND2X1 AND_tmp153 (.Y(ttmp153),.A(N2129),.B(N1171));
AND2X1 AND_tmp154 (.Y(ttmp154),.A(N2286),.B(ttmp153));
AND2X1 AND_tmp155 (.Y(ttmp155),.A(N2427),.B(ttmp154));
AND2X1 AND_tmp156 (.Y(N2639),.A(N2361),.B(ttmp155));
AND2X1 AND_tmp157 (.Y(ttmp157),.A(N2119),.B(N1171));
AND2X1 AND_tmp158 (.Y(ttmp158),.A(N2297),.B(ttmp157));
AND2X1 AND_tmp159 (.Y(ttmp159),.A(N2427),.B(ttmp158));
AND2X1 AND_tmp160 (.Y(N2642),.A(N2361),.B(ttmp159));
AND2X1 AND_tmp161 (.Y(ttmp161),.A(N2104),.B(N1171));
AND2X1 AND_tmp162 (.Y(ttmp162),.A(N2297),.B(ttmp161));
AND2X1 AND_tmp163 (.Y(ttmp163),.A(N2427),.B(ttmp162));
AND2X1 AND_tmp164 (.Y(N2645),.A(N2375),.B(ttmp163));
AND2X1 AND_tmp165 (.Y(ttmp165),.A(N2143),.B(N1171));
AND2X1 AND_tmp166 (.Y(ttmp166),.A(N2297),.B(ttmp165));
AND2X1 AND_tmp167 (.Y(ttmp167),.A(N2427),.B(ttmp166));
AND2X1 AND_tmp168 (.Y(N2648),.A(N2340),.B(ttmp167));
AND2X1 AND_tmp169 (.Y(ttmp169),.A(N2129),.B(N1188));
AND2X1 AND_tmp170 (.Y(ttmp170),.A(N2297),.B(ttmp169));
AND2X1 AND_tmp171 (.Y(ttmp171),.A(N2427),.B(ttmp170));
AND2X1 AND_tmp172 (.Y(N2651),.A(N2353),.B(ttmp171));
AND2X1 AND_tmp173 (.Y(ttmp173),.A(N2129),.B(N1188));
AND2X1 AND_tmp174 (.Y(ttmp174),.A(N2386),.B(ttmp173));
AND2X1 AND_tmp175 (.Y(ttmp175),.A(N2326),.B(ttmp174));
AND2X1 AND_tmp176 (.Y(N2655),.A(N2361),.B(ttmp175));
AND2X1 AND_tmp177 (.Y(ttmp177),.A(N2119),.B(N1188));
AND2X1 AND_tmp178 (.Y(ttmp178),.A(N2386),.B(ttmp177));
AND2X1 AND_tmp179 (.Y(ttmp179),.A(N2326),.B(ttmp178));
AND2X1 AND_tmp180 (.Y(N2658),.A(N2361),.B(ttmp179));
AND2X1 AND_tmp181 (.Y(ttmp181),.A(N2104),.B(N1188));
AND2X1 AND_tmp182 (.Y(ttmp182),.A(N2386),.B(ttmp181));
AND2X1 AND_tmp183 (.Y(ttmp183),.A(N2326),.B(ttmp182));
AND2X1 AND_tmp184 (.Y(N2661),.A(N2375),.B(ttmp183));
AND2X1 AND_tmp185 (.Y(ttmp185),.A(N2129),.B(N1188));
AND2X1 AND_tmp186 (.Y(ttmp186),.A(N2386),.B(ttmp185));
AND2X1 AND_tmp187 (.Y(ttmp187),.A(N2326),.B(ttmp186));
AND2X1 AND_tmp188 (.Y(N2664),.A(N2353),.B(ttmp187));
NAND2X1 NAND2_750 (.Y(N2669),.A(N2558),.B(N534));
INVX1 NOT1_751 (.Y(N2670),.A(N2558));
NAND2X1 NAND2_752 (.Y(N2671),.A(N2561),.B(N535));
INVX1 NOT1_753 (.Y(N2672),.A(N2561));
NAND2X1 NAND2_754 (.Y(N2673),.A(N2564),.B(N536));
INVX1 NOT1_755 (.Y(N2674),.A(N2564));
NAND2X1 NAND2_756 (.Y(N2675),.A(N2567),.B(N537));
INVX1 NOT1_757 (.Y(N2676),.A(N2567));
NAND2X1 NAND2_758 (.Y(N2682),.A(N2570),.B(N543));
INVX1 NOT1_759 (.Y(N2683),.A(N2570));
NAND2X1 NAND2_760 (.Y(N2688),.A(N2573),.B(N548));
INVX1 NOT1_761 (.Y(N2689),.A(N2573));
NAND2X1 NAND2_762 (.Y(N2690),.A(N2576),.B(N549));
INVX1 NOT1_763 (.Y(N2691),.A(N2576));
AND2X1 AND_tmp189 (.Y(ttmp189),.A(N2633),.B(N2634));
AND2X1 AND_tmp190 (.Y(ttmp190),.A(N2627),.B(ttmp189));
AND2X1 AND_tmp191 (.Y(ttmp191),.A(N2628),.B(ttmp190));
AND2X1 AND_tmp192 (.Y(ttmp192),.A(N2629),.B(ttmp191));
AND2X1 AND_tmp193 (.Y(ttmp193),.A(N2630),.B(ttmp192));
AND2X1 AND_tmp194 (.Y(ttmp194),.A(N2631),.B(ttmp193));
AND2X1 AND_tmp195 (.Y(N2710),.A(N2632),.B(ttmp194));
NAND2X1 NAND2_765 (.Y(N2720),.A(N343),.B(N2670));
NAND2X1 NAND2_766 (.Y(N2721),.A(N346),.B(N2672));
NAND2X1 NAND2_767 (.Y(N2722),.A(N349),.B(N2674));
NAND2X1 NAND2_768 (.Y(N2723),.A(N352),.B(N2676));
NAND2X1 NAND2_769 (.Y(N2724),.A(N2639),.B(N538));
INVX1 NOT1_770 (.Y(N2725),.A(N2639));
NAND2X1 NAND2_771 (.Y(N2726),.A(N2642),.B(N539));
INVX1 NOT1_772 (.Y(N2727),.A(N2642));
NAND2X1 NAND2_773 (.Y(N2728),.A(N2645),.B(N540));
INVX1 NOT1_774 (.Y(N2729),.A(N2645));
NAND2X1 NAND2_775 (.Y(N2730),.A(N2648),.B(N541));
INVX1 NOT1_776 (.Y(N2731),.A(N2648));
NAND2X1 NAND2_777 (.Y(N2732),.A(N2651),.B(N542));
INVX1 NOT1_778 (.Y(N2733),.A(N2651));
NAND2X1 NAND2_779 (.Y(N2734),.A(N370),.B(N2683));
NAND2X1 NAND2_780 (.Y(N2735),.A(N2655),.B(N544));
INVX1 NOT1_781 (.Y(N2736),.A(N2655));
NAND2X1 NAND2_782 (.Y(N2737),.A(N2658),.B(N545));
INVX1 NOT1_783 (.Y(N2738),.A(N2658));
NAND2X1 NAND2_784 (.Y(N2739),.A(N2661),.B(N546));
INVX1 NOT1_785 (.Y(N2740),.A(N2661));
NAND2X1 NAND2_786 (.Y(N2741),.A(N2664),.B(N547));
INVX1 NOT1_787 (.Y(N2742),.A(N2664));
NAND2X1 NAND2_788 (.Y(N2743),.A(N385),.B(N2689));
NAND2X1 NAND2_789 (.Y(N2744),.A(N388),.B(N2691));
AND2X1 AND_tmp196 (.Y(ttmp196),.A(N2600),.B(N2603));
AND2X1 AND_tmp197 (.Y(ttmp197),.A(N2537),.B(ttmp196));
AND2X1 AND_tmp198 (.Y(ttmp198),.A(N2540),.B(ttmp197));
AND2X1 AND_tmp199 (.Y(ttmp199),.A(N2543),.B(ttmp198));
AND2X1 AND_tmp200 (.Y(ttmp200),.A(N2546),.B(ttmp199));
AND2X1 AND_tmp201 (.Y(ttmp201),.A(N2594),.B(ttmp200));
NAND2X1 NAND_tmp202 (.Y(N2745),.A(N2597),.B(ttmp201));
AND2X1 AND_tmp203 (.Y(ttmp203),.A(N2552),.B(N2555));
AND2X1 AND_tmp204 (.Y(ttmp204),.A(N2606),.B(ttmp203));
AND2X1 AND_tmp205 (.Y(ttmp205),.A(N2549),.B(ttmp204));
AND2X1 AND_tmp206 (.Y(ttmp206),.A(N2611),.B(ttmp205));
AND2X1 AND_tmp207 (.Y(ttmp207),.A(N2614),.B(ttmp206));
AND2X1 AND_tmp208 (.Y(ttmp208),.A(N2617),.B(ttmp207));
NAND2X1 NAND_tmp209 (.Y(N2746),.A(N2620),.B(ttmp208));
AND2X1 AND_tmp210 (.Y(ttmp210),.A(N2600),.B(N2603));
AND2X1 AND_tmp211 (.Y(ttmp211),.A(N2537),.B(ttmp210));
AND2X1 AND_tmp212 (.Y(ttmp212),.A(N2540),.B(ttmp211));
AND2X1 AND_tmp213 (.Y(ttmp213),.A(N2543),.B(ttmp212));
AND2X1 AND_tmp214 (.Y(ttmp214),.A(N2546),.B(ttmp213));
AND2X1 AND_tmp215 (.Y(ttmp215),.A(N2594),.B(ttmp214));
AND2X1 AND_tmp216 (.Y(N2747),.A(N2597),.B(ttmp215));
AND2X1 AND_tmp217 (.Y(ttmp217),.A(N2552),.B(N2555));
AND2X1 AND_tmp218 (.Y(ttmp218),.A(N2606),.B(ttmp217));
AND2X1 AND_tmp219 (.Y(ttmp219),.A(N2549),.B(ttmp218));
AND2X1 AND_tmp220 (.Y(ttmp220),.A(N2611),.B(ttmp219));
AND2X1 AND_tmp221 (.Y(ttmp221),.A(N2614),.B(ttmp220));
AND2X1 AND_tmp222 (.Y(ttmp222),.A(N2617),.B(ttmp221));
AND2X1 AND_tmp223 (.Y(N2750),.A(N2620),.B(ttmp222));
NAND2X1 NAND2_794 (.Y(N2753),.A(N2669),.B(N2720));
NAND2X1 NAND2_795 (.Y(N2754),.A(N2671),.B(N2721));
NAND2X1 NAND2_796 (.Y(N2755),.A(N2673),.B(N2722));
NAND2X1 NAND2_797 (.Y(N2756),.A(N2675),.B(N2723));
NAND2X1 NAND2_798 (.Y(N2757),.A(N355),.B(N2725));
NAND2X1 NAND2_799 (.Y(N2758),.A(N358),.B(N2727));
NAND2X1 NAND2_800 (.Y(N2759),.A(N361),.B(N2729));
NAND2X1 NAND2_801 (.Y(N2760),.A(N364),.B(N2731));
NAND2X1 NAND2_802 (.Y(N2761),.A(N367),.B(N2733));
NAND2X1 NAND2_803 (.Y(N2762),.A(N2682),.B(N2734));
NAND2X1 NAND2_804 (.Y(N2763),.A(N373),.B(N2736));
NAND2X1 NAND2_805 (.Y(N2764),.A(N376),.B(N2738));
NAND2X1 NAND2_806 (.Y(N2765),.A(N379),.B(N2740));
NAND2X1 NAND2_807 (.Y(N2766),.A(N382),.B(N2742));
NAND2X1 NAND2_808 (.Y(N2767),.A(N2688),.B(N2743));
NAND2X1 NAND2_809 (.Y(N2768),.A(N2690),.B(N2744));
AND2X1 AND2_810 (.Y(N2773),.A(N2745),.B(N275));
AND2X1 AND2_811 (.Y(N2776),.A(N2746),.B(N276));
NAND2X1 NAND2_812 (.Y(N2779),.A(N2724),.B(N2757));
NAND2X1 NAND2_813 (.Y(N2780),.A(N2726),.B(N2758));
NAND2X1 NAND2_814 (.Y(N2781),.A(N2728),.B(N2759));
NAND2X1 NAND2_815 (.Y(N2782),.A(N2730),.B(N2760));
NAND2X1 NAND2_816 (.Y(N2783),.A(N2732),.B(N2761));
NAND2X1 NAND2_817 (.Y(N2784),.A(N2735),.B(N2763));
NAND2X1 NAND2_818 (.Y(N2785),.A(N2737),.B(N2764));
NAND2X1 NAND2_819 (.Y(N2786),.A(N2739),.B(N2765));
NAND2X1 NAND2_820 (.Y(N2787),.A(N2741),.B(N2766));
AND2X1 AND_tmp224 (.Y(ttmp224),.A(N2750),.B(N2710));
AND2X1 AND_tmp225 (.Y(N2788),.A(N2747),.B(ttmp224));
NAND2X1 NAND2_822 (.Y(N2789),.A(N2747),.B(N2750));
AND2X1 AND_tmp226 (.Y(ttmp226),.A(N99),.B(N2788));
AND2X1 AND_tmp227 (.Y(ttmp227),.A(N338),.B(ttmp226));
AND2X1 AND_tmp228 (.Y(N2800),.A(N2279),.B(ttmp227));
NAND2X1 NAND2_824 (.Y(N2807),.A(N2773),.B(N2018));
INVX1 NOT1_825 (.Y(N2808),.A(N2773));
NAND2X1 NAND2_826 (.Y(N2809),.A(N2776),.B(N2019));
INVX1 NOT1_827 (.Y(N2810),.A(N2776));
NOR2X1 NOR2_828 (.Y(N2811),.A(N2384),.B(N2800));
AND2X1 AND_tmp229 (.Y(ttmp229),.A(N283),.B(N2789));
AND2X1 AND_tmp230 (.Y(N2812),.A(N897),.B(ttmp229));
AND2X1 AND_tmp231 (.Y(ttmp231),.A(N283),.B(N2789));
AND2X1 AND_tmp232 (.Y(N2815),.A(N76),.B(ttmp231));
AND2X1 AND_tmp233 (.Y(ttmp233),.A(N283),.B(N2789));
AND2X1 AND_tmp234 (.Y(N2818),.A(N82),.B(ttmp233));
AND2X1 AND_tmp235 (.Y(ttmp235),.A(N283),.B(N2789));
AND2X1 AND_tmp236 (.Y(N2821),.A(N85),.B(ttmp235));
AND2X1 AND_tmp237 (.Y(ttmp237),.A(N283),.B(N2789));
AND2X1 AND_tmp238 (.Y(N2824),.A(N898),.B(ttmp237));
NAND2X1 NAND2_834 (.Y(N2827),.A(N1965),.B(N2808));
NAND2X1 NAND2_835 (.Y(N2828),.A(N1968),.B(N2810));
AND2X1 AND_tmp239 (.Y(ttmp239),.A(N283),.B(N2789));
AND2X1 AND_tmp240 (.Y(N2829),.A(N79),.B(ttmp239));
NAND2X1 NAND2_837 (.Y(N2843),.A(N2807),.B(N2827));
NAND2X1 NAND2_838 (.Y(N2846),.A(N2809),.B(N2828));
NAND2X1 NAND2_839 (.Y(N2850),.A(N2812),.B(N2076));
NAND2X1 NAND2_840 (.Y(N2851),.A(N2815),.B(N2077));
NAND2X1 NAND2_841 (.Y(N2852),.A(N2818),.B(N1915));
NAND2X1 NAND2_842 (.Y(N2853),.A(N2821),.B(N1857));
NAND2X1 NAND2_843 (.Y(N2854),.A(N2824),.B(N1938));
INVX1 NOT1_844 (.Y(N2857),.A(N2812));
INVX1 NOT1_845 (.Y(N2858),.A(N2815));
INVX1 NOT1_846 (.Y(N2859),.A(N2818));
INVX1 NOT1_847 (.Y(N2860),.A(N2821));
INVX1 NOT1_848 (.Y(N2861),.A(N2824));
INVX1 NOT1_849 (.Y(N2862),.A(N2829));
NAND2X1 NAND2_850 (.Y(N2863),.A(N2829),.B(N1985));
NAND2X1 NAND2_851 (.Y(N2866),.A(N2052),.B(N2857));
NAND2X1 NAND2_852 (.Y(N2867),.A(N2055),.B(N2858));
NAND2X1 NAND2_853 (.Y(N2868),.A(N1866),.B(N2859));
NAND2X1 NAND2_854 (.Y(N2869),.A(N1818),.B(N2860));
NAND2X1 NAND2_855 (.Y(N2870),.A(N1902),.B(N2861));
NAND2X1 NAND2_856 (.Y(N2871),.A(N2843),.B(N886));
INVX1 NOT1_857 (.Y(N2872),.A(N2843));
NAND2X1 NAND2_858 (.Y(N2873),.A(N2846),.B(N887));
INVX1 NOT1_859 (.Y(N2874),.A(N2846));
NAND2X1 NAND2_860 (.Y(N2875),.A(N1933),.B(N2862));
NAND2X1 NAND2_861 (.Y(N2876),.A(N2866),.B(N2850));
NAND2X1 NAND2_862 (.Y(N2877),.A(N2867),.B(N2851));
NAND2X1 NAND2_863 (.Y(N2878),.A(N2868),.B(N2852));
NAND2X1 NAND2_864 (.Y(N2879),.A(N2869),.B(N2853));
NAND2X1 NAND2_865 (.Y(N2880),.A(N2870),.B(N2854));
NAND2X1 NAND2_866 (.Y(N2881),.A(N682),.B(N2872));
NAND2X1 NAND2_867 (.Y(N2882),.A(N685),.B(N2874));
NAND2X1 NAND2_868 (.Y(N2883),.A(N2875),.B(N2863));
AND2X1 AND2_869 (.Y(N2886),.A(N2876),.B(N550));
AND2X1 AND2_870 (.Y(N2887),.A(N551),.B(N2877));
AND2X1 AND2_871 (.Y(N2888),.A(N553),.B(N2878));
AND2X1 AND2_872 (.Y(N2889),.A(N2879),.B(N554));
AND2X1 AND2_873 (.Y(N2890),.A(N555),.B(N2880));
NAND2X1 NAND2_874 (.Y(N2891),.A(N2871),.B(N2881));
NAND2X1 NAND2_875 (.Y(N2892),.A(N2873),.B(N2882));
NAND2X1 NAND2_876 (.Y(N2895),.A(N2883),.B(N1461));
INVX1 NOT1_877 (.Y(N2896),.A(N2883));
NAND2X1 NAND2_878 (.Y(N2897),.A(N1383),.B(N2896));
NAND2X1 NAND2_879 (.Y(N2898),.A(N2895),.B(N2897));
AND2X1 AND2_880 (.Y(N2899),.A(N2898),.B(N552));
endmodule