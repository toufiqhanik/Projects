module c5315 (N1,N4,N11,N14,N17,N20,N23,N24,N25,N26,N27,N31,N34,N37,N40,N43,N46,N49,N52,N53,N54,N61,N64,N67,N70,N73,N76,N79,N80,N81,N82,N83,N86,N87,N88,N91,N94,N97,N100,N103,N106,N109,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N126,N127,N128,N129,N130,N131,N132,N135,N136,N137,N140,N141,N145,N146,N149,N152,N155,N158,N161,N164,N167,N170,N173,N176,N179,N182,N185,N188,N191,N194,N197,N200,N203,N206,N209,N210,N217,N218,N225,N226,N233,N234,N241,N242,N245,N248,N251,N254,N257,N264,N265,N272,N273,N280,N281,N288,N289,N292,N293,N299,N302,N307,N308,N315,N316,N323,N324,N331,N332,N335,N338,N341,N348,N351,N358,N361,N366,N369,N372,N373,N374,N386,N389,N400,N411,N422,N435,N446,N457,N468,N479,N490,N503,N514,N523,N534,N545,N549,N552,N556,N559,N562,N566,N571,N574,N577,N580,N583,N588,N591,N592,N595,N596,N597,N598,N599,N603,N607,N610,N613,N616,N619,N625,N631,N709,N816,N1066,N1137,N1138,N1139,N1140,N1141,N1142,N1143,N1144,N1145,N1147,N1152,N1153,N1154,N1155,N1972,N2054,N2060,N2061,N2139,N2142,N2309,N2387,N2527,N2584,N2590,N2623,N3357,N3358,N3359,N3360,N3604,N3613,N4272,N4275,N4278,N4279,N4737,N4738,N4739,N4740,N5240,N5388,N6641,N6643,N6646,N6648,N6716,N6877,N6924,N6925,N6926,N6927,N7015,N7363,N7365,N7432,N7449,N7465,N7466,N7467,N7469,N7470,N7471,N7472,N7473,N7474,N7476,N7503,N7504,N7506,N7511,N7515,N7516,N7517,N7518,N7519,N7520,N7521,N7522,N7600,N7601,N7602,N7603,N7604,N7605,N7606,N7607,N7626,N7698,N7699,N7700,N7701,N7702,N7703,N7704,N7705,N7706,N7707,N7735,N7736,N7737,N7738,N7739,N7740,N7741,N7742,N7754,N7755,N7756,N7757,N7758,N7759,N7760,N7761,N8075,N8076,N8123,N8124,N8127,N8128,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11);
input N1,N4,N11,N14,N17,N20,N23,N24,N25,N26,N27,N31,N34,N37,N40,N43,N46,N49,N52,N53,N54,N61,N64,N67,N70,N73,N76,N79,N80,N81,N82,N83,N86,N87,N88,N91,N94,N97,N100,N103,N106,N109,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N126,N127,N128,N129,N130,N131,N132,N135,N136,N137,N140,N141,N145,N146,N149,N152,N155,N158,N161,N164,N167,N170,N173,N176,N179,N182,N185,N188,N191,N194,N197,N200,N203,N206,N209,N210,N217,N218,N225,N226,N233,N234,N241,N242,N245,N248,N251,N254,N257,N264,N265,N272,N273,N280,N281,N288,N289,N292,N293,N299,N302,N307,N308,N315,N316,N323,N324,N331,N332,N335,N338,N341,N348,N351,N358,N361,N366,N369,N372,N373,N374,N386,N389,N400,N411,N422,N435,N446,N457,N468,N479,N490,N503,N514,N523,N534,N545,N549,N552,N556,N559,N562,N566,N571,N574,N577,N580,N583,N588,N591,N592,N595,N596,N597,N598,N599,N603,N607,N610,N613,N616,N619,N625,N631,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11;
output N709,N816,N1066,N1137,N1138,N1139,N1140,N1141,N1142,N1143,N1144,N1145,N1147,N1152,N1153,N1154,N1155,N1972,N2054,N2060,N2061,N2139,N2142,N2309,N2387,N2527,N2584,N2590,N2623,N3357,N3358,N3359,N3360,N3604,N3613,N4272,N4275,N4278,N4279,N4737,N4738,N4739,N4740,N5240,N5388,N6641,N6643,N6646,N6648,N6716,N6877,N6924,N6925,N6926,N6927,N7015,N7363,N7365,N7432,N7449,N7465,N7466,N7467,N7469,N7470,N7471,N7472,N7473,N7474,N7476,N7503,N7504,N7506,N7511,N7515,N7516,N7517,N7518,N7519,N7520,N7521,N7522,N7600,N7601,N7602,N7603,N7604,N7605,N7606,N7607,N7626,N7698,N7699,N7700,N7701,N7702,N7703,N7704,N7705,N7706,N7707,N7735,N7736,N7737,N7738,N7739,N7740,N7741,N7742,N7754,N7755,N7756,N7757,N7758,N7759,N7760,N7761,N8075,N8076,N8123,N8124,N8127,N8128;
wire N1042,N1043,N1067,N1080,N1092,N1104,N1146,N1148,N1149,N1150,N1151,N1156,N1157,N1161,N1173,N1185,N1197,N1209,N1213,N1216,N1219,N1223,N1235,N1247,N1259,N1271,N1280,N1292,N1303,N1315,N1327,N1339,N1351,N1363,N1375,N1378,N1381,N1384,N1387,N1390,N1393,N1396,N1415,N1418,N1421,N1424,N1427,N1430,N1433,N1436,N1455,N1462,N1469,N1475,N1479,N1482,N1492,N1495,N1498,N1501,N1504,N1507,N1510,N1513,N1516,N1519,N1522,N1525,N1542,N1545,N1548,N1551,N1554,N1557,N1560,N1563,N1566,N1573,N1580,N1583,N1588,N1594,N1597,N1600,N1603,N1606,N1609,N1612,N1615,N1618,N1621,N1624,N1627,N1630,N1633,N1636,N1639,N1642,N1645,N1648,N1651,N1654,N1657,N1660,N1663,N1675,N1685,N1697,N1709,N1721,N1727,N1731,N1743,N1755,N1758,N1761,N1769,N1777,N1785,N1793,N1800,N1807,N1814,N1821,N1824,N1827,N1830,N1833,N1836,N1839,N1842,N1845,N1848,N1851,N1854,N1857,N1860,N1863,N1866,N1869,N1872,N1875,N1878,N1881,N1884,N1887,N1890,N1893,N1896,N1899,N1902,N1905,N1908,N1911,N1914,N1917,N1920,N1923,N1926,N1929,N1932,N1935,N1938,N1941,N1944,N1947,N1950,N1953,N1956,N1959,N1962,N1965,N1968,N2349,N2350,N2585,N2586,N2587,N2588,N2589,N2591,N2592,N2593,N2594,N2595,N2596,N2597,N2598,N2599,N2600,N2601,N2602,N2603,N2604,N2605,N2606,N2607,N2608,N2609,N2610,N2611,N2612,N2613,N2614,N2615,N2616,N2617,N2618,N2619,N2620,N2621,N2622,N2624,N2625,N2626,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,N2635,N2636,N2637,N2638,N2639,N2640,N2641,N2642,N2643,N2644,N2645,N2646,N2647,N2653,N2664,N2675,N2681,N2692,N2703,N2704,N2709,N2710,N2711,N2712,N2713,N2714,N2715,N2716,N2717,N2718,N2719,N2720,N2721,N2722,N2728,N2739,N2750,N2756,N2767,N2778,N2779,N2790,N2801,N2812,N2823,N2824,N2825,N2826,N2827,N2828,N2829,N2830,N2831,N2832,N2833,N2834,N2835,N2836,N2837,N2838,N2839,N2840,N2841,N2842,N2843,N2844,N2845,N2846,N2847,N2848,N2849,N2850,N2851,N2852,N2853,N2854,N2855,N2861,N2867,N2868,N2869,N2870,N2871,N2872,N2873,N2874,N2875,N2876,N2877,N2882,N2891,N2901,N2902,N2903,N2904,N2905,N2906,N2907,N2908,N2909,N2910,N2911,N2912,N2913,N2914,N2915,N2916,N2917,N2918,N2919,N2920,N2921,N2922,N2923,N2924,N2925,N2926,N2927,N2928,N2929,N2930,N2931,N2932,N2933,N2934,N2935,N2936,N2937,N2938,N2939,N2940,N2941,N2942,N2948,N2954,N2955,N2956,N2957,N2958,N2959,N2960,N2961,N2962,N2963,N2964,N2969,N2970,N2971,N2972,N2973,N2974,N2975,N2976,N2977,N2978,N2979,N2980,N2981,N2982,N2983,N2984,N2985,N2986,N2987,N2988,N2989,N2990,N2991,N2992,N2993,N2994,N2995,N2996,N2997,N2998,N2999,N3000,N3003,N3006,N3007,N3010,N3013,N3014,N3015,N3016,N3017,N3018,N3019,N3020,N3021,N3022,N3023,N3024,N3025,N3026,N3027,N3028,N3029,N3030,N3031,N3032,N3033,N3034,N3035,N3038,N3041,N3052,N3063,N3068,N3071,N3072,N3073,N3074,N3075,N3086,N3097,N3108,N3119,N3130,N3141,N3142,N3143,N3144,N3145,N3146,N3147,N3158,N3169,N3180,N3191,N3194,N3195,N3196,N3197,N3198,N3199,N3200,N3203,N3401,N3402,N3403,N3404,N3405,N3406,N3407,N3408,N3409,N3410,N3411,N3412,N3413,N3414,N3415,N3416,N3444,N3445,N3446,N3447,N3448,N3449,N3450,N3451,N3452,N3453,N3454,N3455,N3456,N3459,N3460,N3461,N3462,N3463,N3464,N3465,N3466,N3481,N3482,N3483,N3484,N3485,N3486,N3487,N3488,N3489,N3490,N3491,N3492,N3493,N3502,N3503,N3504,N3505,N3506,N3507,N3508,N3509,N3510,N3511,N3512,N3513,N3514,N3515,N3558,N3559,N3560,N3561,N3562,N3563,N3605,N3606,N3607,N3608,N3609,N3610,N3614,N3615,N3616,N3617,N3618,N3619,N3620,N3621,N3622,N3623,N3624,N3625,N3626,N3627,N3628,N3629,N3630,N3631,N3632,N3633,N3634,N3635,N3636,N3637,N3638,N3639,N3640,N3641,N3642,N3643,N3644,N3645,N3646,N3647,N3648,N3649,N3650,N3651,N3652,N3653,N3654,N3655,N3656,N3657,N3658,N3659,N3660,N3661,N3662,N3663,N3664,N3665,N3666,N3667,N3668,N3669,N3670,N3671,N3672,N3673,N3674,N3675,N3676,N3677,N3678,N3679,N3680,N3681,N3682,N3683,N3684,N3685,N3686,N3687,N3688,N3689,N3691,N3700,N3701,N3702,N3703,N3704,N3705,N3708,N3709,N3710,N3711,N3712,N3713,N3715,N3716,N3717,N3718,N3719,N3720,N3721,N3722,N3723,N3724,N3725,N3726,N3727,N3728,N3729,N3730,N3731,N3732,N3738,N3739,N3740,N3741,N3742,N3743,N3744,N3745,N3746,N3747,N3748,N3749,N3750,N3751,N3752,N3753,N3754,N3755,N3756,N3757,N3758,N3759,N3760,N3761,N3762,N3763,N3764,N3765,N3766,N3767,N3768,N3769,N3770,N3771,N3775,N3779,N3780,N3781,N3782,N3783,N3784,N3785,N3786,N3787,N3788,N3789,N3793,N3797,N3800,N3801,N3802,N3803,N3804,N3805,N3806,N3807,N3808,N3809,N3810,N3813,N3816,N3819,N3822,N3823,N3824,N3827,N3828,N3829,N3830,N3831,N3834,N3835,N3836,N3837,N3838,N3839,N3840,N3841,N3842,N3849,N3855,N3861,N3867,N3873,N3881,N3887,N3893,N3908,N3909,N3911,N3914,N3915,N3916,N3917,N3918,N3919,N3920,N3921,N3927,N3933,N3942,N3948,N3956,N3962,N3968,N3975,N3976,N3977,N3978,N3979,N3980,N3981,N3982,N3983,N3984,N3987,N3988,N3989,N3990,N3991,N3998,N4008,N4011,N4021,N4024,N4027,N4031,N4032,N4033,N4034,N4035,N4036,N4037,N4038,N4039,N4040,N4041,N4042,N4067,N4080,N4088,N4091,N4094,N4097,N4100,N4103,N4106,N4109,N4144,N4147,N4150,N4153,N4156,N4159,N4183,N4184,N4185,N4186,N4188,N4191,N4196,N4197,N4198,N4199,N4200,N4203,N4206,N4209,N4212,N4215,N4219,N4223,N4224,N4225,N4228,N4231,N4234,N4237,N4240,N4243,N4246,N4249,N4252,N4255,N4258,N4263,N4264,N4267,N4268,N4269,N4270,N4271,N4273,N4274,N4276,N4277,N4280,N4284,N4290,N4297,N4298,N4301,N4305,N4310,N4316,N4320,N4325,N4331,N4332,N4336,N4342,N4349,N4357,N4364,N4375,N4379,N4385,N4392,N4396,N4400,N4405,N4412,N4418,N4425,N4436,N4440,N4445,N4451,N4456,N4462,N4469,N4477,N4512,N4515,N4516,N4521,N4523,N4524,N4532,N4547,N4548,N4551,N4554,N4557,N4560,N4563,N4566,N4569,N4572,N4575,N4578,N4581,N4584,N4587,N4590,N4593,N4596,N4599,N4602,N4605,N4608,N4611,N4614,N4617,N4621,N4624,N4627,N4630,N4633,N4637,N4640,N4643,N4646,N4649,N4652,N4655,N4658,N4662,N4665,N4668,N4671,N4674,N4677,N4680,N4683,N4686,N4689,N4692,N4695,N4698,N4701,N4702,N4720,N4721,N4724,N4725,N4726,N4727,N4728,N4729,N4730,N4731,N4732,N4733,N4734,N4735,N4736,N4741,N4855,N4856,N4908,N4909,N4939,N4942,N4947,N4953,N4954,N4955,N4956,N4957,N4958,N4959,N4960,N4961,N4965,N4966,N4967,N4968,N4972,N4973,N4974,N4975,N4976,N4977,N4978,N4979,N4980,N4981,N4982,N4983,N4984,N4985,N4986,N4987,N5049,N5052,N5053,N5054,N5055,N5056,N5057,N5058,N5059,N5060,N5061,N5062,N5063,N5065,N5066,N5067,N5068,N5069,N5070,N5071,N5072,N5073,N5074,N5075,N5076,N5077,N5078,N5079,N5080,N5081,N5082,N5083,N5084,N5085,N5086,N5087,N5088,N5089,N5090,N5091,N5092,N5093,N5094,N5095,N5096,N5097,N5098,N5099,N5100,N5101,N5102,N5103,N5104,N5105,N5106,N5107,N5108,N5109,N5110,N5111,N5112,N5113,N5114,N5115,N5116,N5117,N5118,N5119,N5120,N5121,N5122,N5123,N5124,N5125,N5126,N5127,N5128,N5129,N5130,N5131,N5132,N5133,N5135,N5136,N5137,N5138,N5139,N5140,N5141,N5142,N5143,N5144,N5145,N5146,N5147,N5148,N5150,N5153,N5154,N5155,N5156,N5157,N5160,N5161,N5162,N5163,N5164,N5165,N5166,N5169,N5172,N5173,N5176,N5177,N5180,N5183,N5186,N5189,N5192,N5195,N5198,N5199,N5202,N5205,N5208,N5211,N5214,N5217,N5220,N5223,N5224,N5225,N5226,N5227,N5228,N5229,N5230,N5232,N5233,N5234,N5235,N5236,N5239,N5241,N5242,N5243,N5244,N5245,N5246,N5247,N5248,N5249,N5250,N5252,N5253,N5254,N5255,N5256,N5257,N5258,N5259,N5260,N5261,N5262,N5263,N5264,N5274,N5275,N5282,N5283,N5284,N5298,N5299,N5300,N5303,N5304,N5305,N5306,N5307,N5308,N5309,N5310,N5311,N5312,N5315,N5319,N5324,N5328,N5331,N5332,N5346,N5363,N5364,N5365,N5366,N5367,N5368,N5369,N5370,N5371,N5374,N5377,N5382,N5385,N5389,N5396,N5407,N5418,N5424,N5431,N5441,N5452,N5462,N5469,N5470,N5477,N5488,N5498,N5506,N5520,N5536,N5549,N5555,N5562,N5573,N5579,N5595,N5606,N5616,N5617,N5618,N5619,N5620,N5621,N5622,N5624,N5634,N5655,N5671,N5684,N5690,N5691,N5692,N5696,N5700,N5703,N5707,N5711,N5726,N5727,N5728,N5730,N5731,N5732,N5733,N5734,N5735,N5736,N5739,N5742,N5745,N5755,N5756,N5954,N5955,N5956,N6005,N6006,N6023,N6024,N6025,N6028,N6031,N6034,N6037,N6040,N6044,N6045,N6048,N6051,N6054,N6065,N6066,N6067,N6068,N6069,N6071,N6072,N6073,N6074,N6075,N6076,N6077,N6078,N6079,N6080,N6083,N6084,N6085,N6086,N6087,N6088,N6089,N6090,N6091,N6094,N6095,N6096,N6097,N6098,N6099,N6100,N6101,N6102,N6103,N6104,N6105,N6106,N6107,N6108,N6111,N6112,N6113,N6114,N6115,N6116,N6117,N6120,N6121,N6122,N6123,N6124,N6125,N6126,N6127,N6128,N6129,N6130,N6131,N6132,N6133,N6134,N6135,N6136,N6137,N6138,N6139,N6140,N6143,N6144,N6145,N6146,N6147,N6148,N6149,N6152,N6153,N6154,N6155,N6156,N6157,N6158,N6159,N6160,N6161,N6162,N6163,N6164,N6168,N6171,N6172,N6173,N6174,N6175,N6178,N6179,N6180,N6181,N6182,N6183,N6184,N6185,N6186,N6187,N6188,N6189,N6190,N6191,N6192,N6193,N6194,N6197,N6200,N6203,N6206,N6209,N6212,N6215,N6218,N6221,N6234,N6235,N6238,N6241,N6244,N6247,N6250,N6253,N6256,N6259,N6262,N6265,N6268,N6271,N6274,N6277,N6280,N6283,N6286,N6289,N6292,N6295,N6298,N6301,N6304,N6307,N6310,N6313,N6316,N6319,N6322,N6325,N6328,N6331,N6335,N6338,N6341,N6344,N6347,N6350,N6353,N6356,N6359,N6364,N6367,N6370,N6373,N6374,N6375,N6376,N6377,N6378,N6382,N6386,N6388,N6392,N6397,N6411,N6415,N6419,N6427,N6434,N6437,N6441,N6445,N6448,N6449,N6466,N6469,N6470,N6471,N6472,N6473,N6474,N6475,N6476,N6477,N6478,N6482,N6486,N6490,N6494,N6500,N6504,N6508,N6512,N6516,N6526,N6536,N6539,N6553,N6556,N6566,N6569,N6572,N6575,N6580,N6584,N6587,N6592,N6599,N6606,N6609,N6619,N6622,N6630,N6631,N6632,N6633,N6634,N6637,N6640,N6650,N6651,N6653,N6655,N6657,N6659,N6660,N6661,N6662,N6663,N6664,N6666,N6668,N6670,N6672,N6675,N6680,N6681,N6682,N6683,N6689,N6690,N6691,N6692,N6693,N6695,N6698,N6699,N6700,N6703,N6708,N6709,N6710,N6711,N6712,N6713,N6714,N6715,N6718,N6719,N6720,N6721,N6722,N6724,N6739,N6740,N6741,N6744,N6745,N6746,N6751,N6752,N6753,N6754,N6755,N6760,N6761,N6762,N6772,N6773,N6776,N6777,N6782,N6783,N6784,N6785,N6790,N6791,N6792,N6795,N6801,N6802,N6803,N6804,N6805,N6806,N6807,N6808,N6809,N6810,N6811,N6812,N6813,N6814,N6815,N6816,N6817,N6823,N6824,N6825,N6826,N6827,N6828,N6829,N6830,N6831,N6834,N6835,N6836,N6837,N6838,N6839,N6840,N6841,N6842,N6843,N6844,N6850,N6851,N6852,N6853,N6854,N6855,N6856,N6857,N6860,N6861,N6862,N6863,N6866,N6872,N6873,N6874,N6875,N6876,N6879,N6880,N6881,N6884,N6885,N6888,N6889,N6890,N6891,N6894,N6895,N6896,N6897,N6900,N6901,N6904,N6905,N6908,N6909,N6912,N6913,N6914,N6915,N6916,N6919,N6922,N6923,N6930,N6932,N6935,N6936,N6937,N6938,N6939,N6940,N6946,N6947,N6948,N6949,N6953,N6954,N6955,N6956,N6957,N6958,N6964,N6965,N6966,N6967,N6973,N6974,N6975,N6976,N6977,N6978,N6979,N6987,N6990,N6999,N7002,N7003,N7006,N7011,N7012,N7013,N7016,N7018,N7019,N7020,N7021,N7022,N7023,N7028,N7031,N7034,N7037,N7040,N7041,N7044,N7045,N7046,N7047,N7048,N7049,N7054,N7057,N7060,N7064,N7065,N7072,N7073,N7074,N7075,N7076,N7079,N7080,N7083,N7084,N7085,N7086,N7087,N7088,N7089,N7090,N7093,N7094,N7097,N7101,N7105,N7110,N7114,N7115,N7116,N7125,N7126,N7127,N7130,N7131,N7139,N7140,N7141,N7146,N7147,N7149,N7150,N7151,N7152,N7153,N7158,N7159,N7160,N7166,N7167,N7168,N7169,N7170,N7171,N7172,N7173,N7174,N7175,N7176,N7177,N7178,N7179,N7180,N7181,N7182,N7183,N7184,N7185,N7186,N7187,N7188,N7189,N7190,N7196,N7197,N7198,N7204,N7205,N7206,N7207,N7208,N7209,N7212,N7215,N7216,N7217,N7218,N7219,N7222,N7225,N7228,N7229,N7236,N7239,N7242,N7245,N7250,N7257,N7260,N7263,N7268,N7269,N7270,N7276,N7282,N7288,N7294,N7300,N7301,N7304,N7310,N7320,N7321,N7328,N7338,N7339,N7340,N7341,N7342,N7349,N7357,N7364,N7394,N7397,N7402,N7405,N7406,N7407,N7408,N7409,N7412,N7415,N7416,N7417,N7418,N7419,N7420,N7421,N7424,N7425,N7426,N7427,N7428,N7429,N7430,N7431,N7433,N7434,N7435,N7436,N7437,N7438,N7439,N7440,N7441,N7442,N7443,N7444,N7445,N7446,N7447,N7448,N7450,N7451,N7452,N7453,N7454,N7455,N7456,N7457,N7458,N7459,N7460,N7461,N7462,N7463,N7464,N7468,N7479,N7481,N7482,N7483,N7484,N7485,N7486,N7487,N7488,N7489,N7492,N7493,N7498,N7499,N7500,N7505,N7507,N7508,N7509,N7510,N7512,N7513,N7514,N7525,N7526,N7527,N7528,N7529,N7530,N7531,N7537,N7543,N7549,N7555,N7561,N7567,N7573,N7579,N7582,N7585,N7586,N7587,N7588,N7589,N7592,N7595,N7598,N7599,N7624,N7625,N7631,N7636,N7657,N7658,N7665,N7666,N7667,N7668,N7669,N7670,N7671,N7672,N7673,N7674,N7675,N7676,N7677,N7678,N7679,N7680,N7681,N7682,N7683,N7684,N7685,N7686,N7687,N7688,N7689,N7690,N7691,N7692,N7693,N7694,N7695,N7696,N7697,N7708,N7709,N7710,N7711,N7712,N7715,N7718,N7719,N7720,N7721,N7722,N7723,N7724,N7727,N7728,N7729,N7730,N7731,N7732,N7733,N7734,N7743,N7744,N7749,N7750,N7751,N7762,N7765,N7768,N7769,N7770,N7771,N7772,N7775,N7778,N7781,N7782,N7787,N7788,N7795,N7796,N7797,N7798,N7799,N7800,N7803,N7806,N7807,N7808,N7809,N7810,N7811,N7812,N7815,N7816,N7821,N7822,N7823,N7826,N7829,N7832,N7833,N7834,N7835,N7836,N7839,N7842,N7845,N7846,N7851,N7852,N7859,N7860,N7861,N7862,N7863,N7864,N7867,N7870,N7871,N7872,N7873,N7874,N7875,N7876,N7879,N7880,N7885,N7886,N7887,N7890,N7893,N7896,N7897,N7898,N7899,N7900,N7903,N7906,N7909,N7910,N7917,N7918,N7923,N7924,N7925,N7926,N7927,N7928,N7929,N7930,N7931,N7932,N7935,N7938,N7939,N7940,N7943,N7944,N7945,N7946,N7951,N7954,N7957,N7960,N7963,N7966,N7967,N7968,N7969,N7970,N7973,N7974,N7984,N7985,N7987,N7988,N7989,N7990,N7991,N7992,N7993,N7994,N7995,N7996,N7997,N7998,N8001,N8004,N8009,N8013,N8017,N8020,N8021,N8022,N8023,N8025,N8026,N8027,N8031,N8032,N8033,N8034,N8035,N8036,N8037,N8038,N8039,N8040,N8041,N8042,N8043,N8044,N8045,N8048,N8055,N8056,N8057,N8058,N8059,N8060,N8061,N8064,N8071,N8072,N8073,N8074,N8077,N8078,N8079,N8082,N8089,N8090,N8091,N8092,N8093,N8096,N8099,N8102,N8113,N8114,N8115,N8116,N8117,N8118,N8119,N8120,N8121,N8122,N8125,N8126,compare0,compare1,compare2,compare3,compare4,compare5,compare6,compare7,compare8,compare9,compare10,compare11,andgate0,andgate1,andgate2,andgate3,andgate4,andgate5,andgate6,andgate7,andgate8,andgate9,andgate10,orgate0,orgate1,orgate2,orgate3,orgate4,orgate5,orgate6,orgate7,orgate8,orgate9,orgate10,andgate11,N709_sar;
BUFX1 BUFF1_1 (.Y(N709_sar),.A(N141));
BUFX1 BUFF1_2 (.Y(N816),.A(N293));
AND2X1 AND2_3 (.Y(N1042),.A(N135),.B(N631));
INVX1 NOT1_4 (.Y(N1043),.A(N591));
BUFX1 BUFF1_5 (.Y(N1066),.A(N592));
INVX1 NOT1_6 (.Y(N1067),.A(N595));
INVX1 NOT1_7 (.Y(N1080),.A(N596));
INVX1 NOT1_8 (.Y(N1092),.A(N597));
INVX1 NOT1_9 (.Y(N1104),.A(N598));
INVX1 NOT1_10 (.Y(N1137),.A(N545));
INVX1 NOT1_11 (.Y(N1138),.A(N348));
INVX1 NOT1_12 (.Y(N1139),.A(N366));
AND2X1 AND2_13 (.Y(N1140),.A(N552),.B(N562));
INVX1 NOT1_14 (.Y(N1141),.A(N549));
INVX1 NOT1_15 (.Y(N1142),.A(N545));
INVX1 NOT1_16 (.Y(N1143),.A(N545));
INVX1 NOT1_17 (.Y(N1144),.A(N338));
INVX1 NOT1_18 (.Y(N1145),.A(N358));
NAND2X1 NAND2_19 (.Y(N1146),.A(N373),.B(N1));
AND2X1 AND2_20 (.Y(N1147),.A(N141),.B(N145));
INVX1 NOT1_21 (.Y(N1148),.A(N592));
INVX1 NOT1_22 (.Y(N1149),.A(N1042));
AND2X1 AND2_23 (.Y(N1150),.A(N1043),.B(N27));
AND2X1 AND2_24 (.Y(N1151),.A(N386),.B(N556));
INVX1 NOT1_25 (.Y(N1152),.A(N245));
INVX1 NOT1_26 (.Y(N1153),.A(N552));
INVX1 NOT1_27 (.Y(N1154),.A(N562));
INVX1 NOT1_28 (.Y(N1155),.A(N559));
AND2X1 AND_tmp1 (.Y(ttmp1),.A(N556),.B(N552));
AND2X1 AND_tmp2 (.Y(ttmp2),.A(N386),.B(ttmp1));
AND2X1 AND_tmp3 (.Y(N1156),.A(N559),.B(ttmp2));
INVX1 NOT1_30 (.Y(N1157),.A(N566));
BUFX1 BUFF1_31 (.Y(N1161),.A(N571));
BUFX1 BUFF1_32 (.Y(N1173),.A(N574));
BUFX1 BUFF1_33 (.Y(N1185),.A(N571));
BUFX1 BUFF1_34 (.Y(N1197),.A(N574));
BUFX1 BUFF1_35 (.Y(N1209),.A(N137));
BUFX1 BUFF1_36 (.Y(N1213),.A(N137));
BUFX1 BUFF1_37 (.Y(N1216),.A(N141));
INVX1 NOT1_38 (.Y(N1219),.A(N583));
BUFX1 BUFF1_39 (.Y(N1223),.A(N577));
BUFX1 BUFF1_40 (.Y(N1235),.A(N580));
BUFX1 BUFF1_41 (.Y(N1247),.A(N577));
BUFX1 BUFF1_42 (.Y(N1259),.A(N580));
BUFX1 BUFF1_43 (.Y(N1271),.A(N254));
BUFX1 BUFF1_44 (.Y(N1280),.A(N251));
BUFX1 BUFF1_45 (.Y(N1292),.A(N251));
BUFX1 BUFF1_46 (.Y(N1303),.A(N248));
BUFX1 BUFF1_47 (.Y(N1315),.A(N248));
BUFX1 BUFF1_48 (.Y(N1327),.A(N610));
BUFX1 BUFF1_49 (.Y(N1339),.A(N607));
BUFX1 BUFF1_50 (.Y(N1351),.A(N613));
BUFX1 BUFF1_51 (.Y(N1363),.A(N616));
BUFX1 BUFF1_52 (.Y(N1375),.A(N210));
BUFX1 BUFF1_53 (.Y(N1378),.A(N210));
BUFX1 BUFF1_54 (.Y(N1381),.A(N218));
BUFX1 BUFF1_55 (.Y(N1384),.A(N218));
BUFX1 BUFF1_56 (.Y(N1387),.A(N226));
BUFX1 BUFF1_57 (.Y(N1390),.A(N226));
BUFX1 BUFF1_58 (.Y(N1393),.A(N234));
BUFX1 BUFF1_59 (.Y(N1396),.A(N234));
BUFX1 BUFF1_60 (.Y(N1415),.A(N257));
BUFX1 BUFF1_61 (.Y(N1418),.A(N257));
BUFX1 BUFF1_62 (.Y(N1421),.A(N265));
BUFX1 BUFF1_63 (.Y(N1424),.A(N265));
BUFX1 BUFF1_64 (.Y(N1427),.A(N273));
BUFX1 BUFF1_65 (.Y(N1430),.A(N273));
BUFX1 BUFF1_66 (.Y(N1433),.A(N281));
BUFX1 BUFF1_67 (.Y(N1436),.A(N281));
BUFX1 BUFF1_68 (.Y(N1455),.A(N335));
BUFX1 BUFF1_69 (.Y(N1462),.A(N335));
BUFX1 BUFF1_70 (.Y(N1469),.A(N206));
AND2X1 AND2_71 (.Y(N1475),.A(N27),.B(N31));
BUFX1 BUFF1_72 (.Y(N1479),.A(N1));
BUFX1 BUFF1_73 (.Y(N1482),.A(N588));
BUFX1 BUFF1_74 (.Y(N1492),.A(N293));
BUFX1 BUFF1_75 (.Y(N1495),.A(N302));
BUFX1 BUFF1_76 (.Y(N1498),.A(N308));
BUFX1 BUFF1_77 (.Y(N1501),.A(N308));
BUFX1 BUFF1_78 (.Y(N1504),.A(N316));
BUFX1 BUFF1_79 (.Y(N1507),.A(N316));
BUFX1 BUFF1_80 (.Y(N1510),.A(N324));
BUFX1 BUFF1_81 (.Y(N1513),.A(N324));
BUFX1 BUFF1_82 (.Y(N1516),.A(N341));
BUFX1 BUFF1_83 (.Y(N1519),.A(N341));
BUFX1 BUFF1_84 (.Y(N1522),.A(N351));
BUFX1 BUFF1_85 (.Y(N1525),.A(N351));
BUFX1 BUFF1_86 (.Y(N1542),.A(N257));
BUFX1 BUFF1_87 (.Y(N1545),.A(N257));
BUFX1 BUFF1_88 (.Y(N1548),.A(N265));
BUFX1 BUFF1_89 (.Y(N1551),.A(N265));
BUFX1 BUFF1_90 (.Y(N1554),.A(N273));
BUFX1 BUFF1_91 (.Y(N1557),.A(N273));
BUFX1 BUFF1_92 (.Y(N1560),.A(N281));
BUFX1 BUFF1_93 (.Y(N1563),.A(N281));
BUFX1 BUFF1_94 (.Y(N1566),.A(N332));
BUFX1 BUFF1_95 (.Y(N1573),.A(N332));
BUFX1 BUFF1_96 (.Y(N1580),.A(N549));
AND2X1 AND2_97 (.Y(N1583),.A(N31),.B(N27));
INVX1 NOT1_98 (.Y(N1588),.A(N588));
BUFX1 BUFF1_99 (.Y(N1594),.A(N324));
BUFX1 BUFF1_100 (.Y(N1597),.A(N324));
BUFX1 BUFF1_101 (.Y(N1600),.A(N341));
BUFX1 BUFF1_102 (.Y(N1603),.A(N341));
BUFX1 BUFF1_103 (.Y(N1606),.A(N351));
BUFX1 BUFF1_104 (.Y(N1609),.A(N351));
BUFX1 BUFF1_105 (.Y(N1612),.A(N293));
BUFX1 BUFF1_106 (.Y(N1615),.A(N302));
BUFX1 BUFF1_107 (.Y(N1618),.A(N308));
BUFX1 BUFF1_108 (.Y(N1621),.A(N308));
BUFX1 BUFF1_109 (.Y(N1624),.A(N316));
BUFX1 BUFF1_110 (.Y(N1627),.A(N316));
BUFX1 BUFF1_111 (.Y(N1630),.A(N361));
BUFX1 BUFF1_112 (.Y(N1633),.A(N361));
BUFX1 BUFF1_113 (.Y(N1636),.A(N210));
BUFX1 BUFF1_114 (.Y(N1639),.A(N210));
BUFX1 BUFF1_115 (.Y(N1642),.A(N218));
BUFX1 BUFF1_116 (.Y(N1645),.A(N218));
BUFX1 BUFF1_117 (.Y(N1648),.A(N226));
BUFX1 BUFF1_118 (.Y(N1651),.A(N226));
BUFX1 BUFF1_119 (.Y(N1654),.A(N234));
BUFX1 BUFF1_120 (.Y(N1657),.A(N234));
INVX1 NOT1_121 (.Y(N1660),.A(N324));
BUFX1 BUFF1_122 (.Y(N1663),.A(N242));
BUFX1 BUFF1_123 (.Y(N1675),.A(N242));
BUFX1 BUFF1_124 (.Y(N1685),.A(N254));
BUFX1 BUFF1_125 (.Y(N1697),.A(N610));
BUFX1 BUFF1_126 (.Y(N1709),.A(N607));
BUFX1 BUFF1_127 (.Y(N1721),.A(N625));
BUFX1 BUFF1_128 (.Y(N1727),.A(N619));
BUFX1 BUFF1_129 (.Y(N1731),.A(N613));
BUFX1 BUFF1_130 (.Y(N1743),.A(N616));
INVX1 NOT1_131 (.Y(N1755),.A(N599));
INVX1 NOT1_132 (.Y(N1758),.A(N603));
BUFX1 BUFF1_133 (.Y(N1761),.A(N619));
BUFX1 BUFF1_134 (.Y(N1769),.A(N625));
BUFX1 BUFF1_135 (.Y(N1777),.A(N619));
BUFX1 BUFF1_136 (.Y(N1785),.A(N625));
BUFX1 BUFF1_137 (.Y(N1793),.A(N619));
BUFX1 BUFF1_138 (.Y(N1800),.A(N625));
BUFX1 BUFF1_139 (.Y(N1807),.A(N619));
BUFX1 BUFF1_140 (.Y(N1814),.A(N625));
BUFX1 BUFF1_141 (.Y(N1821),.A(N299));
BUFX1 BUFF1_142 (.Y(N1824),.A(N446));
BUFX1 BUFF1_143 (.Y(N1827),.A(N457));
BUFX1 BUFF1_144 (.Y(N1830),.A(N468));
BUFX1 BUFF1_145 (.Y(N1833),.A(N422));
BUFX1 BUFF1_146 (.Y(N1836),.A(N435));
BUFX1 BUFF1_147 (.Y(N1839),.A(N389));
BUFX1 BUFF1_148 (.Y(N1842),.A(N400));
BUFX1 BUFF1_149 (.Y(N1845),.A(N411));
BUFX1 BUFF1_150 (.Y(N1848),.A(N374));
BUFX1 BUFF1_151 (.Y(N1851),.A(N4));
BUFX1 BUFF1_152 (.Y(N1854),.A(N446));
BUFX1 BUFF1_153 (.Y(N1857),.A(N457));
BUFX1 BUFF1_154 (.Y(N1860),.A(N468));
BUFX1 BUFF1_155 (.Y(N1863),.A(N435));
BUFX1 BUFF1_156 (.Y(N1866),.A(N389));
BUFX1 BUFF1_157 (.Y(N1869),.A(N400));
BUFX1 BUFF1_158 (.Y(N1872),.A(N411));
BUFX1 BUFF1_159 (.Y(N1875),.A(N422));
BUFX1 BUFF1_160 (.Y(N1878),.A(N374));
BUFX1 BUFF1_161 (.Y(N1881),.A(N479));
BUFX1 BUFF1_162 (.Y(N1884),.A(N490));
BUFX1 BUFF1_163 (.Y(N1887),.A(N503));
BUFX1 BUFF1_164 (.Y(N1890),.A(N514));
BUFX1 BUFF1_165 (.Y(N1893),.A(N523));
BUFX1 BUFF1_166 (.Y(N1896),.A(N534));
BUFX1 BUFF1_167 (.Y(N1899),.A(N54));
BUFX1 BUFF1_168 (.Y(N1902),.A(N479));
BUFX1 BUFF1_169 (.Y(N1905),.A(N503));
BUFX1 BUFF1_170 (.Y(N1908),.A(N514));
BUFX1 BUFF1_171 (.Y(N1911),.A(N523));
BUFX1 BUFF1_172 (.Y(N1914),.A(N534));
BUFX1 BUFF1_173 (.Y(N1917),.A(N490));
BUFX1 BUFF1_174 (.Y(N1920),.A(N361));
BUFX1 BUFF1_175 (.Y(N1923),.A(N369));
BUFX1 BUFF1_176 (.Y(N1926),.A(N341));
BUFX1 BUFF1_177 (.Y(N1929),.A(N351));
BUFX1 BUFF1_178 (.Y(N1932),.A(N308));
BUFX1 BUFF1_179 (.Y(N1935),.A(N316));
BUFX1 BUFF1_180 (.Y(N1938),.A(N293));
BUFX1 BUFF1_181 (.Y(N1941),.A(N302));
BUFX1 BUFF1_182 (.Y(N1944),.A(N281));
BUFX1 BUFF1_183 (.Y(N1947),.A(N289));
BUFX1 BUFF1_184 (.Y(N1950),.A(N265));
BUFX1 BUFF1_185 (.Y(N1953),.A(N273));
BUFX1 BUFF1_186 (.Y(N1956),.A(N234));
BUFX1 BUFF1_187 (.Y(N1959),.A(N257));
BUFX1 BUFF1_188 (.Y(N1962),.A(N218));
BUFX1 BUFF1_189 (.Y(N1965),.A(N226));
BUFX1 BUFF1_190 (.Y(N1968),.A(N210));
INVX1 NOT1_191 (.Y(N1972),.A(N1146));
AND2X1 AND2_192 (.Y(N2054),.A(N136),.B(N1148));
INVX1 NOT1_193 (.Y(N2060),.A(N1150));
INVX1 NOT1_194 (.Y(N2061),.A(N1151));
BUFX1 BUFF1_195 (.Y(N2139),.A(N1209));
BUFX1 BUFF1_196 (.Y(N2142),.A(N1216));
BUFX1 BUFF1_197 (.Y(N2309),.A(N1479));
AND2X1 AND2_198 (.Y(N2349),.A(N1104),.B(N514));
OR2X1 OR2_199 (.Y(N2350),.A(N1067),.B(N514));
BUFX1 BUFF1_200 (.Y(N2387),.A(N1580));
BUFX1 BUFF1_201 (.Y(N2527),.A(N1821));
INVX1 NOT1_202 (.Y(N2584),.A(N1580));
AND2X1 AND_tmp4 (.Y(ttmp4),.A(N1161),.B(N1173));
AND2X1 AND_tmp5 (.Y(N2585),.A(N170),.B(ttmp4));
AND2X1 AND_tmp6 (.Y(ttmp6),.A(N1161),.B(N1173));
AND2X1 AND_tmp7 (.Y(N2586),.A(N173),.B(ttmp6));
AND2X1 AND_tmp8 (.Y(ttmp8),.A(N1161),.B(N1173));
AND2X1 AND_tmp9 (.Y(N2587),.A(N167),.B(ttmp8));
AND2X1 AND_tmp10 (.Y(ttmp10),.A(N1161),.B(N1173));
AND2X1 AND_tmp11 (.Y(N2588),.A(N164),.B(ttmp10));
AND2X1 AND_tmp12 (.Y(ttmp12),.A(N1161),.B(N1173));
AND2X1 AND_tmp13 (.Y(N2589),.A(N161),.B(ttmp12));
NAND2X1 NAND2_208 (.Y(N2590),.A(N1475),.B(N140));
AND2X1 AND_tmp14 (.Y(ttmp14),.A(N1185),.B(N1197));
AND2X1 AND_tmp15 (.Y(N2591),.A(N185),.B(ttmp14));
AND2X1 AND_tmp16 (.Y(ttmp16),.A(N1185),.B(N1197));
AND2X1 AND_tmp17 (.Y(N2592),.A(N158),.B(ttmp16));
AND2X1 AND_tmp18 (.Y(ttmp18),.A(N1185),.B(N1197));
AND2X1 AND_tmp19 (.Y(N2593),.A(N152),.B(ttmp18));
AND2X1 AND_tmp20 (.Y(ttmp20),.A(N1185),.B(N1197));
AND2X1 AND_tmp21 (.Y(N2594),.A(N146),.B(ttmp20));
AND2X1 AND_tmp22 (.Y(ttmp22),.A(N1223),.B(N1235));
AND2X1 AND_tmp23 (.Y(N2595),.A(N170),.B(ttmp22));
AND2X1 AND_tmp24 (.Y(ttmp24),.A(N1223),.B(N1235));
AND2X1 AND_tmp25 (.Y(N2596),.A(N173),.B(ttmp24));
AND2X1 AND_tmp26 (.Y(ttmp26),.A(N1223),.B(N1235));
AND2X1 AND_tmp27 (.Y(N2597),.A(N167),.B(ttmp26));
AND2X1 AND_tmp28 (.Y(ttmp28),.A(N1223),.B(N1235));
AND2X1 AND_tmp29 (.Y(N2598),.A(N164),.B(ttmp28));
AND2X1 AND_tmp30 (.Y(ttmp30),.A(N1223),.B(N1235));
AND2X1 AND_tmp31 (.Y(N2599),.A(N161),.B(ttmp30));
AND2X1 AND_tmp32 (.Y(ttmp32),.A(N1247),.B(N1259));
AND2X1 AND_tmp33 (.Y(N2600),.A(N185),.B(ttmp32));
AND2X1 AND_tmp34 (.Y(ttmp34),.A(N1247),.B(N1259));
AND2X1 AND_tmp35 (.Y(N2601),.A(N158),.B(ttmp34));
AND2X1 AND_tmp36 (.Y(ttmp36),.A(N1247),.B(N1259));
AND2X1 AND_tmp37 (.Y(N2602),.A(N152),.B(ttmp36));
AND2X1 AND_tmp38 (.Y(ttmp38),.A(N1247),.B(N1259));
AND2X1 AND_tmp39 (.Y(N2603),.A(N146),.B(ttmp38));
AND2X1 AND_tmp40 (.Y(ttmp40),.A(N1731),.B(N1743));
AND2X1 AND_tmp41 (.Y(N2604),.A(N106),.B(ttmp40));
AND2X1 AND_tmp42 (.Y(ttmp42),.A(N1327),.B(N1339));
AND2X1 AND_tmp43 (.Y(N2605),.A(N61),.B(ttmp42));
AND2X1 AND_tmp44 (.Y(ttmp44),.A(N1697),.B(N1709));
AND2X1 AND_tmp45 (.Y(N2606),.A(N106),.B(ttmp44));
AND2X1 AND_tmp46 (.Y(ttmp46),.A(N1697),.B(N1709));
AND2X1 AND_tmp47 (.Y(N2607),.A(N49),.B(ttmp46));
AND2X1 AND_tmp48 (.Y(ttmp48),.A(N1697),.B(N1709));
AND2X1 AND_tmp49 (.Y(N2608),.A(N103),.B(ttmp48));
AND2X1 AND_tmp50 (.Y(ttmp50),.A(N1697),.B(N1709));
AND2X1 AND_tmp51 (.Y(N2609),.A(N40),.B(ttmp50));
AND2X1 AND_tmp52 (.Y(ttmp52),.A(N1697),.B(N1709));
AND2X1 AND_tmp53 (.Y(N2610),.A(N37),.B(ttmp52));
AND2X1 AND_tmp54 (.Y(ttmp54),.A(N1327),.B(N1339));
AND2X1 AND_tmp55 (.Y(N2611),.A(N20),.B(ttmp54));
AND2X1 AND_tmp56 (.Y(ttmp56),.A(N1327),.B(N1339));
AND2X1 AND_tmp57 (.Y(N2612),.A(N17),.B(ttmp56));
AND2X1 AND_tmp58 (.Y(ttmp58),.A(N1327),.B(N1339));
AND2X1 AND_tmp59 (.Y(N2613),.A(N70),.B(ttmp58));
AND2X1 AND_tmp60 (.Y(ttmp60),.A(N1327),.B(N1339));
AND2X1 AND_tmp61 (.Y(N2614),.A(N64),.B(ttmp60));
AND2X1 AND_tmp62 (.Y(ttmp62),.A(N1731),.B(N1743));
AND2X1 AND_tmp63 (.Y(N2615),.A(N49),.B(ttmp62));
AND2X1 AND_tmp64 (.Y(ttmp64),.A(N1731),.B(N1743));
AND2X1 AND_tmp65 (.Y(N2616),.A(N103),.B(ttmp64));
AND2X1 AND_tmp66 (.Y(ttmp66),.A(N1731),.B(N1743));
AND2X1 AND_tmp67 (.Y(N2617),.A(N40),.B(ttmp66));
AND2X1 AND_tmp68 (.Y(ttmp68),.A(N1731),.B(N1743));
AND2X1 AND_tmp69 (.Y(N2618),.A(N37),.B(ttmp68));
AND2X1 AND_tmp70 (.Y(ttmp70),.A(N1351),.B(N1363));
AND2X1 AND_tmp71 (.Y(N2619),.A(N20),.B(ttmp70));
AND2X1 AND_tmp72 (.Y(ttmp72),.A(N1351),.B(N1363));
AND2X1 AND_tmp73 (.Y(N2620),.A(N17),.B(ttmp72));
AND2X1 AND_tmp74 (.Y(ttmp74),.A(N1351),.B(N1363));
AND2X1 AND_tmp75 (.Y(N2621),.A(N70),.B(ttmp74));
AND2X1 AND_tmp76 (.Y(ttmp76),.A(N1351),.B(N1363));
AND2X1 AND_tmp77 (.Y(N2622),.A(N64),.B(ttmp76));
INVX1 NOT1_241 (.Y(N2623),.A(N1475));
AND2X1 AND_tmp78 (.Y(ttmp78),.A(N1758),.B(N599));
AND2X1 AND_tmp79 (.Y(N2624),.A(N123),.B(ttmp78));
AND2X1 AND2_243 (.Y(N2625),.A(N1777),.B(N1785));
AND2X1 AND_tmp80 (.Y(ttmp80),.A(N1351),.B(N1363));
AND2X1 AND_tmp81 (.Y(N2626),.A(N61),.B(ttmp80));
AND2X1 AND2_245 (.Y(N2627),.A(N1761),.B(N1769));
INVX1 NOT1_246 (.Y(N2628),.A(N1824));
INVX1 NOT1_247 (.Y(N2629),.A(N1827));
INVX1 NOT1_248 (.Y(N2630),.A(N1830));
INVX1 NOT1_249 (.Y(N2631),.A(N1833));
INVX1 NOT1_250 (.Y(N2632),.A(N1836));
INVX1 NOT1_251 (.Y(N2633),.A(N1839));
INVX1 NOT1_252 (.Y(N2634),.A(N1842));
INVX1 NOT1_253 (.Y(N2635),.A(N1845));
INVX1 NOT1_254 (.Y(N2636),.A(N1848));
INVX1 NOT1_255 (.Y(N2637),.A(N1851));
INVX1 NOT1_256 (.Y(N2638),.A(N1854));
INVX1 NOT1_257 (.Y(N2639),.A(N1857));
INVX1 NOT1_258 (.Y(N2640),.A(N1860));
INVX1 NOT1_259 (.Y(N2641),.A(N1863));
INVX1 NOT1_260 (.Y(N2642),.A(N1866));
INVX1 NOT1_261 (.Y(N2643),.A(N1869));
INVX1 NOT1_262 (.Y(N2644),.A(N1872));
INVX1 NOT1_263 (.Y(N2645),.A(N1875));
INVX1 NOT1_264 (.Y(N2646),.A(N1878));
BUFX1 BUFF1_265 (.Y(N2647),.A(N1209));
INVX1 NOT1_266 (.Y(N2653),.A(N1161));
INVX1 NOT1_267 (.Y(N2664),.A(N1173));
BUFX1 BUFF1_268 (.Y(N2675),.A(N1209));
INVX1 NOT1_269 (.Y(N2681),.A(N1185));
INVX1 NOT1_270 (.Y(N2692),.A(N1197));
AND2X1 AND_tmp82 (.Y(ttmp82),.A(N1185),.B(N1197));
AND2X1 AND_tmp83 (.Y(N2703),.A(N179),.B(ttmp82));
BUFX1 BUFF1_272 (.Y(N2704),.A(N1479));
INVX1 NOT1_273 (.Y(N2709),.A(N1881));
INVX1 NOT1_274 (.Y(N2710),.A(N1884));
INVX1 NOT1_275 (.Y(N2711),.A(N1887));
INVX1 NOT1_276 (.Y(N2712),.A(N1890));
INVX1 NOT1_277 (.Y(N2713),.A(N1893));
INVX1 NOT1_278 (.Y(N2714),.A(N1896));
INVX1 NOT1_279 (.Y(N2715),.A(N1899));
INVX1 NOT1_280 (.Y(N2716),.A(N1902));
INVX1 NOT1_281 (.Y(N2717),.A(N1905));
INVX1 NOT1_282 (.Y(N2718),.A(N1908));
INVX1 NOT1_283 (.Y(N2719),.A(N1911));
INVX1 NOT1_284 (.Y(N2720),.A(N1914));
INVX1 NOT1_285 (.Y(N2721),.A(N1917));
BUFX1 BUFF1_286 (.Y(N2722),.A(N1213));
INVX1 NOT1_287 (.Y(N2728),.A(N1223));
INVX1 NOT1_288 (.Y(N2739),.A(N1235));
BUFX1 BUFF1_289 (.Y(N2750),.A(N1213));
INVX1 NOT1_290 (.Y(N2756),.A(N1247));
INVX1 NOT1_291 (.Y(N2767),.A(N1259));
AND2X1 AND_tmp84 (.Y(ttmp84),.A(N1247),.B(N1259));
AND2X1 AND_tmp85 (.Y(N2778),.A(N179),.B(ttmp84));
INVX1 NOT1_293 (.Y(N2779),.A(N1327));
INVX1 NOT1_294 (.Y(N2790),.A(N1339));
INVX1 NOT1_295 (.Y(N2801),.A(N1351));
INVX1 NOT1_296 (.Y(N2812),.A(N1363));
INVX1 NOT1_297 (.Y(N2823),.A(N1375));
INVX1 NOT1_298 (.Y(N2824),.A(N1378));
INVX1 NOT1_299 (.Y(N2825),.A(N1381));
INVX1 NOT1_300 (.Y(N2826),.A(N1384));
INVX1 NOT1_301 (.Y(N2827),.A(N1387));
INVX1 NOT1_302 (.Y(N2828),.A(N1390));
INVX1 NOT1_303 (.Y(N2829),.A(N1393));
INVX1 NOT1_304 (.Y(N2830),.A(N1396));
AND2X1 AND_tmp86 (.Y(ttmp86),.A(N457),.B(N1378));
AND2X1 AND_tmp87 (.Y(N2831),.A(N1104),.B(ttmp86));
AND2X1 AND_tmp88 (.Y(ttmp88),.A(N468),.B(N1384));
AND2X1 AND_tmp89 (.Y(N2832),.A(N1104),.B(ttmp88));
AND2X1 AND_tmp90 (.Y(ttmp90),.A(N422),.B(N1390));
AND2X1 AND_tmp91 (.Y(N2833),.A(N1104),.B(ttmp90));
AND2X1 AND_tmp92 (.Y(ttmp92),.A(N435),.B(N1396));
AND2X1 AND_tmp93 (.Y(N2834),.A(N1104),.B(ttmp92));
AND2X1 AND2_309 (.Y(N2835),.A(N1067),.B(N1375));
AND2X1 AND2_310 (.Y(N2836),.A(N1067),.B(N1381));
AND2X1 AND2_311 (.Y(N2837),.A(N1067),.B(N1387));
AND2X1 AND2_312 (.Y(N2838),.A(N1067),.B(N1393));
INVX1 NOT1_313 (.Y(N2839),.A(N1415));
INVX1 NOT1_314 (.Y(N2840),.A(N1418));
INVX1 NOT1_315 (.Y(N2841),.A(N1421));
INVX1 NOT1_316 (.Y(N2842),.A(N1424));
INVX1 NOT1_317 (.Y(N2843),.A(N1427));
INVX1 NOT1_318 (.Y(N2844),.A(N1430));
INVX1 NOT1_319 (.Y(N2845),.A(N1433));
INVX1 NOT1_320 (.Y(N2846),.A(N1436));
AND2X1 AND_tmp94 (.Y(ttmp94),.A(N389),.B(N1418));
AND2X1 AND_tmp95 (.Y(N2847),.A(N1104),.B(ttmp94));
AND2X1 AND_tmp96 (.Y(ttmp96),.A(N400),.B(N1424));
AND2X1 AND_tmp97 (.Y(N2848),.A(N1104),.B(ttmp96));
AND2X1 AND_tmp98 (.Y(ttmp98),.A(N411),.B(N1430));
AND2X1 AND_tmp99 (.Y(N2849),.A(N1104),.B(ttmp98));
AND2X1 AND_tmp100 (.Y(ttmp100),.A(N374),.B(N1436));
AND2X1 AND_tmp101 (.Y(N2850),.A(N1104),.B(ttmp100));
AND2X1 AND2_325 (.Y(N2851),.A(N1067),.B(N1415));
AND2X1 AND2_326 (.Y(N2852),.A(N1067),.B(N1421));
AND2X1 AND2_327 (.Y(N2853),.A(N1067),.B(N1427));
AND2X1 AND2_328 (.Y(N2854),.A(N1067),.B(N1433));
INVX1 NOT1_329 (.Y(N2855),.A(N1455));
INVX1 NOT1_330 (.Y(N2861),.A(N1462));
AND2X1 AND2_331 (.Y(N2867),.A(N292),.B(N1455));
AND2X1 AND2_332 (.Y(N2868),.A(N288),.B(N1455));
AND2X1 AND2_333 (.Y(N2869),.A(N280),.B(N1455));
AND2X1 AND2_334 (.Y(N2870),.A(N272),.B(N1455));
AND2X1 AND2_335 (.Y(N2871),.A(N264),.B(N1455));
AND2X1 AND2_336 (.Y(N2872),.A(N241),.B(N1462));
AND2X1 AND2_337 (.Y(N2873),.A(N233),.B(N1462));
AND2X1 AND2_338 (.Y(N2874),.A(N225),.B(N1462));
AND2X1 AND2_339 (.Y(N2875),.A(N217),.B(N1462));
AND2X1 AND2_340 (.Y(N2876),.A(N209),.B(N1462));
BUFX1 BUFF1_341 (.Y(N2877),.A(N1216));
INVX1 NOT1_342 (.Y(N2882),.A(N1482));
INVX1 NOT1_343 (.Y(N2891),.A(N1475));
INVX1 NOT1_344 (.Y(N2901),.A(N1492));
INVX1 NOT1_345 (.Y(N2902),.A(N1495));
INVX1 NOT1_346 (.Y(N2903),.A(N1498));
INVX1 NOT1_347 (.Y(N2904),.A(N1501));
INVX1 NOT1_348 (.Y(N2905),.A(N1504));
INVX1 NOT1_349 (.Y(N2906),.A(N1507));
AND2X1 AND2_350 (.Y(N2907),.A(N1303),.B(N1495));
AND2X1 AND_tmp102 (.Y(ttmp102),.A(N479),.B(N1501));
AND2X1 AND_tmp103 (.Y(N2908),.A(N1303),.B(ttmp102));
AND2X1 AND_tmp104 (.Y(ttmp104),.A(N490),.B(N1507));
AND2X1 AND_tmp105 (.Y(N2909),.A(N1303),.B(ttmp104));
AND2X1 AND2_353 (.Y(N2910),.A(N1663),.B(N1492));
AND2X1 AND2_354 (.Y(N2911),.A(N1663),.B(N1498));
AND2X1 AND2_355 (.Y(N2912),.A(N1663),.B(N1504));
INVX1 NOT1_356 (.Y(N2913),.A(N1510));
INVX1 NOT1_357 (.Y(N2914),.A(N1513));
INVX1 NOT1_358 (.Y(N2915),.A(N1516));
INVX1 NOT1_359 (.Y(N2916),.A(N1519));
INVX1 NOT1_360 (.Y(N2917),.A(N1522));
INVX1 NOT1_361 (.Y(N2918),.A(N1525));
AND2X1 AND_tmp106 (.Y(ttmp106),.A(N503),.B(N1513));
AND2X1 AND_tmp107 (.Y(N2919),.A(N1104),.B(ttmp106));
INVX1 NOT1_363 (.Y(N2920),.A(N2349));
AND2X1 AND_tmp108 (.Y(ttmp108),.A(N523),.B(N1519));
AND2X1 AND_tmp109 (.Y(N2921),.A(N1104),.B(ttmp108));
AND2X1 AND_tmp110 (.Y(ttmp110),.A(N534),.B(N1525));
AND2X1 AND_tmp111 (.Y(N2922),.A(N1104),.B(ttmp110));
AND2X1 AND2_366 (.Y(N2923),.A(N1067),.B(N1510));
AND2X1 AND2_367 (.Y(N2924),.A(N1067),.B(N1516));
AND2X1 AND2_368 (.Y(N2925),.A(N1067),.B(N1522));
INVX1 NOT1_369 (.Y(N2926),.A(N1542));
INVX1 NOT1_370 (.Y(N2927),.A(N1545));
INVX1 NOT1_371 (.Y(N2928),.A(N1548));
INVX1 NOT1_372 (.Y(N2929),.A(N1551));
INVX1 NOT1_373 (.Y(N2930),.A(N1554));
INVX1 NOT1_374 (.Y(N2931),.A(N1557));
INVX1 NOT1_375 (.Y(N2932),.A(N1560));
INVX1 NOT1_376 (.Y(N2933),.A(N1563));
AND2X1 AND_tmp112 (.Y(ttmp112),.A(N389),.B(N1545));
AND2X1 AND_tmp113 (.Y(N2934),.A(N1303),.B(ttmp112));
AND2X1 AND_tmp114 (.Y(ttmp114),.A(N400),.B(N1551));
AND2X1 AND_tmp115 (.Y(N2935),.A(N1303),.B(ttmp114));
AND2X1 AND_tmp116 (.Y(ttmp116),.A(N411),.B(N1557));
AND2X1 AND_tmp117 (.Y(N2936),.A(N1303),.B(ttmp116));
AND2X1 AND_tmp118 (.Y(ttmp118),.A(N374),.B(N1563));
AND2X1 AND_tmp119 (.Y(N2937),.A(N1303),.B(ttmp118));
AND2X1 AND2_381 (.Y(N2938),.A(N1663),.B(N1542));
AND2X1 AND2_382 (.Y(N2939),.A(N1663),.B(N1548));
AND2X1 AND2_383 (.Y(N2940),.A(N1663),.B(N1554));
AND2X1 AND2_384 (.Y(N2941),.A(N1663),.B(N1560));
INVX1 NOT1_385 (.Y(N2942),.A(N1566));
INVX1 NOT1_386 (.Y(N2948),.A(N1573));
AND2X1 AND2_387 (.Y(N2954),.A(N372),.B(N1566));
AND2X1 AND2_388 (.Y(N2955),.A(N366),.B(N1566));
AND2X1 AND2_389 (.Y(N2956),.A(N358),.B(N1566));
AND2X1 AND2_390 (.Y(N2957),.A(N348),.B(N1566));
AND2X1 AND2_391 (.Y(N2958),.A(N338),.B(N1566));
AND2X1 AND2_392 (.Y(N2959),.A(N331),.B(N1573));
AND2X1 AND2_393 (.Y(N2960),.A(N323),.B(N1573));
AND2X1 AND2_394 (.Y(N2961),.A(N315),.B(N1573));
AND2X1 AND2_395 (.Y(N2962),.A(N307),.B(N1573));
AND2X1 AND2_396 (.Y(N2963),.A(N299),.B(N1573));
INVX1 NOT1_397 (.Y(N2964),.A(N1588));
AND2X1 AND2_398 (.Y(N2969),.A(N83),.B(N1588));
AND2X1 AND2_399 (.Y(N2970),.A(N86),.B(N1588));
AND2X1 AND2_400 (.Y(N2971),.A(N88),.B(N1588));
AND2X1 AND2_401 (.Y(N2972),.A(N88),.B(N1588));
INVX1 NOT1_402 (.Y(N2973),.A(N1594));
INVX1 NOT1_403 (.Y(N2974),.A(N1597));
INVX1 NOT1_404 (.Y(N2975),.A(N1600));
INVX1 NOT1_405 (.Y(N2976),.A(N1603));
INVX1 NOT1_406 (.Y(N2977),.A(N1606));
INVX1 NOT1_407 (.Y(N2978),.A(N1609));
AND2X1 AND_tmp120 (.Y(ttmp120),.A(N503),.B(N1597));
AND2X1 AND_tmp121 (.Y(N2979),.A(N1315),.B(ttmp120));
AND2X1 AND2_409 (.Y(N2980),.A(N1315),.B(N514));
AND2X1 AND_tmp122 (.Y(ttmp122),.A(N523),.B(N1603));
AND2X1 AND_tmp123 (.Y(N2981),.A(N1315),.B(ttmp122));
AND2X1 AND_tmp124 (.Y(ttmp124),.A(N534),.B(N1609));
AND2X1 AND_tmp125 (.Y(N2982),.A(N1315),.B(ttmp124));
AND2X1 AND2_412 (.Y(N2983),.A(N1675),.B(N1594));
OR2X1 OR2_413 (.Y(N2984),.A(N1675),.B(N514));
AND2X1 AND2_414 (.Y(N2985),.A(N1675),.B(N1600));
AND2X1 AND2_415 (.Y(N2986),.A(N1675),.B(N1606));
INVX1 NOT1_416 (.Y(N2987),.A(N1612));
INVX1 NOT1_417 (.Y(N2988),.A(N1615));
INVX1 NOT1_418 (.Y(N2989),.A(N1618));
INVX1 NOT1_419 (.Y(N2990),.A(N1621));
INVX1 NOT1_420 (.Y(N2991),.A(N1624));
INVX1 NOT1_421 (.Y(N2992),.A(N1627));
AND2X1 AND2_422 (.Y(N2993),.A(N1315),.B(N1615));
AND2X1 AND_tmp126 (.Y(ttmp126),.A(N479),.B(N1621));
AND2X1 AND_tmp127 (.Y(N2994),.A(N1315),.B(ttmp126));
AND2X1 AND_tmp128 (.Y(ttmp128),.A(N490),.B(N1627));
AND2X1 AND_tmp129 (.Y(N2995),.A(N1315),.B(ttmp128));
AND2X1 AND2_425 (.Y(N2996),.A(N1675),.B(N1612));
AND2X1 AND2_426 (.Y(N2997),.A(N1675),.B(N1618));
AND2X1 AND2_427 (.Y(N2998),.A(N1675),.B(N1624));
INVX1 NOT1_428 (.Y(N2999),.A(N1630));
BUFX1 BUFF1_429 (.Y(N3000),.A(N1469));
BUFX1 BUFF1_430 (.Y(N3003),.A(N1469));
INVX1 NOT1_431 (.Y(N3006),.A(N1633));
BUFX1 BUFF1_432 (.Y(N3007),.A(N1469));
BUFX1 BUFF1_433 (.Y(N3010),.A(N1469));
AND2X1 AND2_434 (.Y(N3013),.A(N1315),.B(N1630));
AND2X1 AND2_435 (.Y(N3014),.A(N1315),.B(N1633));
INVX1 NOT1_436 (.Y(N3015),.A(N1636));
INVX1 NOT1_437 (.Y(N3016),.A(N1639));
INVX1 NOT1_438 (.Y(N3017),.A(N1642));
INVX1 NOT1_439 (.Y(N3018),.A(N1645));
INVX1 NOT1_440 (.Y(N3019),.A(N1648));
INVX1 NOT1_441 (.Y(N3020),.A(N1651));
INVX1 NOT1_442 (.Y(N3021),.A(N1654));
INVX1 NOT1_443 (.Y(N3022),.A(N1657));
AND2X1 AND_tmp130 (.Y(ttmp130),.A(N457),.B(N1639));
AND2X1 AND_tmp131 (.Y(N3023),.A(N1303),.B(ttmp130));
AND2X1 AND_tmp132 (.Y(ttmp132),.A(N468),.B(N1645));
AND2X1 AND_tmp133 (.Y(N3024),.A(N1303),.B(ttmp132));
AND2X1 AND_tmp134 (.Y(ttmp134),.A(N422),.B(N1651));
AND2X1 AND_tmp135 (.Y(N3025),.A(N1303),.B(ttmp134));
AND2X1 AND_tmp136 (.Y(ttmp136),.A(N435),.B(N1657));
AND2X1 AND_tmp137 (.Y(N3026),.A(N1303),.B(ttmp136));
AND2X1 AND2_448 (.Y(N3027),.A(N1663),.B(N1636));
AND2X1 AND2_449 (.Y(N3028),.A(N1663),.B(N1642));
AND2X1 AND2_450 (.Y(N3029),.A(N1663),.B(N1648));
AND2X1 AND2_451 (.Y(N3030),.A(N1663),.B(N1654));
INVX1 NOT1_452 (.Y(N3031),.A(N1920));
INVX1 NOT1_453 (.Y(N3032),.A(N1923));
INVX1 NOT1_454 (.Y(N3033),.A(N1926));
INVX1 NOT1_455 (.Y(N3034),.A(N1929));
BUFX1 BUFF1_456 (.Y(N3035),.A(N1660));
BUFX1 BUFF1_457 (.Y(N3038),.A(N1660));
INVX1 NOT1_458 (.Y(N3041),.A(N1697));
INVX1 NOT1_459 (.Y(N3052),.A(N1709));
INVX1 NOT1_460 (.Y(N3063),.A(N1721));
INVX1 NOT1_461 (.Y(N3068),.A(N1727));
AND2X1 AND2_462 (.Y(N3071),.A(N97),.B(N1721));
AND2X1 AND2_463 (.Y(N3072),.A(N94),.B(N1721));
AND2X1 AND2_464 (.Y(N3073),.A(N97),.B(N1721));
AND2X1 AND2_465 (.Y(N3074),.A(N94),.B(N1721));
INVX1 NOT1_466 (.Y(N3075),.A(N1731));
INVX1 NOT1_467 (.Y(N3086),.A(N1743));
INVX1 NOT1_468 (.Y(N3097),.A(N1761));
INVX1 NOT1_469 (.Y(N3108),.A(N1769));
INVX1 NOT1_470 (.Y(N3119),.A(N1777));
INVX1 NOT1_471 (.Y(N3130),.A(N1785));
INVX1 NOT1_472 (.Y(N3141),.A(N1944));
INVX1 NOT1_473 (.Y(N3142),.A(N1947));
INVX1 NOT1_474 (.Y(N3143),.A(N1950));
INVX1 NOT1_475 (.Y(N3144),.A(N1953));
INVX1 NOT1_476 (.Y(N3145),.A(N1956));
INVX1 NOT1_477 (.Y(N3146),.A(N1959));
INVX1 NOT1_478 (.Y(N3147),.A(N1793));
INVX1 NOT1_479 (.Y(N3158),.A(N1800));
INVX1 NOT1_480 (.Y(N3169),.A(N1807));
INVX1 NOT1_481 (.Y(N3180),.A(N1814));
BUFX1 BUFF1_482 (.Y(N3191),.A(N1821));
INVX1 NOT1_483 (.Y(N3194),.A(N1932));
INVX1 NOT1_484 (.Y(N3195),.A(N1935));
INVX1 NOT1_485 (.Y(N3196),.A(N1938));
INVX1 NOT1_486 (.Y(N3197),.A(N1941));
INVX1 NOT1_487 (.Y(N3198),.A(N1962));
INVX1 NOT1_488 (.Y(N3199),.A(N1965));
BUFX1 BUFF1_489 (.Y(N3200),.A(N1469));
INVX1 NOT1_490 (.Y(N3203),.A(N1968));
BUFX1 BUFF1_491 (.Y(N3357),.A(N2704));
BUFX1 BUFF1_492 (.Y(N3358),.A(N2704));
BUFX1 BUFF1_493 (.Y(N3359),.A(N2704));
BUFX1 BUFF1_494 (.Y(N3360),.A(N2704));
AND2X1 AND_tmp138 (.Y(ttmp138),.A(N1092),.B(N2824));
AND2X1 AND_tmp139 (.Y(N3401),.A(N457),.B(ttmp138));
AND2X1 AND_tmp140 (.Y(ttmp140),.A(N1092),.B(N2826));
AND2X1 AND_tmp141 (.Y(N3402),.A(N468),.B(ttmp140));
AND2X1 AND_tmp142 (.Y(ttmp142),.A(N1092),.B(N2828));
AND2X1 AND_tmp143 (.Y(N3403),.A(N422),.B(ttmp142));
AND2X1 AND_tmp144 (.Y(ttmp144),.A(N1092),.B(N2830));
AND2X1 AND_tmp145 (.Y(N3404),.A(N435),.B(ttmp144));
AND2X1 AND2_499 (.Y(N3405),.A(N1080),.B(N2823));
AND2X1 AND2_500 (.Y(N3406),.A(N1080),.B(N2825));
AND2X1 AND2_501 (.Y(N3407),.A(N1080),.B(N2827));
AND2X1 AND2_502 (.Y(N3408),.A(N1080),.B(N2829));
AND2X1 AND_tmp146 (.Y(ttmp146),.A(N1092),.B(N2840));
AND2X1 AND_tmp147 (.Y(N3409),.A(N389),.B(ttmp146));
AND2X1 AND_tmp148 (.Y(ttmp148),.A(N1092),.B(N2842));
AND2X1 AND_tmp149 (.Y(N3410),.A(N400),.B(ttmp148));
AND2X1 AND_tmp150 (.Y(ttmp150),.A(N1092),.B(N2844));
AND2X1 AND_tmp151 (.Y(N3411),.A(N411),.B(ttmp150));
AND2X1 AND_tmp152 (.Y(ttmp152),.A(N1092),.B(N2846));
AND2X1 AND_tmp153 (.Y(N3412),.A(N374),.B(ttmp152));
AND2X1 AND2_507 (.Y(N3413),.A(N1080),.B(N2839));
AND2X1 AND2_508 (.Y(N3414),.A(N1080),.B(N2841));
AND2X1 AND2_509 (.Y(N3415),.A(N1080),.B(N2843));
AND2X1 AND2_510 (.Y(N3416),.A(N1080),.B(N2845));
AND2X1 AND2_511 (.Y(N3444),.A(N1280),.B(N2902));
AND2X1 AND_tmp154 (.Y(ttmp154),.A(N1280),.B(N2904));
AND2X1 AND_tmp155 (.Y(N3445),.A(N479),.B(ttmp154));
AND2X1 AND_tmp156 (.Y(ttmp156),.A(N1280),.B(N2906));
AND2X1 AND_tmp157 (.Y(N3446),.A(N490),.B(ttmp156));
AND2X1 AND2_514 (.Y(N3447),.A(N1685),.B(N2901));
AND2X1 AND2_515 (.Y(N3448),.A(N1685),.B(N2903));
AND2X1 AND2_516 (.Y(N3449),.A(N1685),.B(N2905));
AND2X1 AND_tmp158 (.Y(ttmp158),.A(N1092),.B(N2914));
AND2X1 AND_tmp159 (.Y(N3450),.A(N503),.B(ttmp158));
AND2X1 AND_tmp160 (.Y(ttmp160),.A(N1092),.B(N2916));
AND2X1 AND_tmp161 (.Y(N3451),.A(N523),.B(ttmp160));
AND2X1 AND_tmp162 (.Y(ttmp162),.A(N1092),.B(N2918));
AND2X1 AND_tmp163 (.Y(N3452),.A(N534),.B(ttmp162));
AND2X1 AND2_520 (.Y(N3453),.A(N1080),.B(N2913));
AND2X1 AND2_521 (.Y(N3454),.A(N1080),.B(N2915));
AND2X1 AND2_522 (.Y(N3455),.A(N1080),.B(N2917));
AND2X1 AND2_523 (.Y(N3456),.A(N2920),.B(N2350));
AND2X1 AND_tmp164 (.Y(ttmp164),.A(N1280),.B(N2927));
AND2X1 AND_tmp165 (.Y(N3459),.A(N389),.B(ttmp164));
AND2X1 AND_tmp166 (.Y(ttmp166),.A(N1280),.B(N2929));
AND2X1 AND_tmp167 (.Y(N3460),.A(N400),.B(ttmp166));
AND2X1 AND_tmp168 (.Y(ttmp168),.A(N1280),.B(N2931));
AND2X1 AND_tmp169 (.Y(N3461),.A(N411),.B(ttmp168));
AND2X1 AND_tmp170 (.Y(ttmp170),.A(N1280),.B(N2933));
AND2X1 AND_tmp171 (.Y(N3462),.A(N374),.B(ttmp170));
AND2X1 AND2_528 (.Y(N3463),.A(N1685),.B(N2926));
AND2X1 AND2_529 (.Y(N3464),.A(N1685),.B(N2928));
AND2X1 AND2_530 (.Y(N3465),.A(N1685),.B(N2930));
AND2X1 AND2_531 (.Y(N3466),.A(N1685),.B(N2932));
AND2X1 AND_tmp172 (.Y(ttmp172),.A(N1292),.B(N2974));
AND2X1 AND_tmp173 (.Y(N3481),.A(N503),.B(ttmp172));
INVX1 NOT1_533 (.Y(N3482),.A(N2980));
AND2X1 AND_tmp174 (.Y(ttmp174),.A(N1292),.B(N2976));
AND2X1 AND_tmp175 (.Y(N3483),.A(N523),.B(ttmp174));
AND2X1 AND_tmp176 (.Y(ttmp176),.A(N1292),.B(N2978));
AND2X1 AND_tmp177 (.Y(N3484),.A(N534),.B(ttmp176));
AND2X1 AND2_536 (.Y(N3485),.A(N1271),.B(N2973));
AND2X1 AND2_537 (.Y(N3486),.A(N1271),.B(N2975));
AND2X1 AND2_538 (.Y(N3487),.A(N1271),.B(N2977));
AND2X1 AND2_539 (.Y(N3488),.A(N1292),.B(N2988));
AND2X1 AND_tmp178 (.Y(ttmp178),.A(N1292),.B(N2990));
AND2X1 AND_tmp179 (.Y(N3489),.A(N479),.B(ttmp178));
AND2X1 AND_tmp180 (.Y(ttmp180),.A(N1292),.B(N2992));
AND2X1 AND_tmp181 (.Y(N3490),.A(N490),.B(ttmp180));
AND2X1 AND2_542 (.Y(N3491),.A(N1271),.B(N2987));
AND2X1 AND2_543 (.Y(N3492),.A(N1271),.B(N2989));
AND2X1 AND2_544 (.Y(N3493),.A(N1271),.B(N2991));
AND2X1 AND2_545 (.Y(N3502),.A(N1292),.B(N2999));
AND2X1 AND2_546 (.Y(N3503),.A(N1292),.B(N3006));
AND2X1 AND_tmp182 (.Y(ttmp182),.A(N1280),.B(N3016));
AND2X1 AND_tmp183 (.Y(N3504),.A(N457),.B(ttmp182));
AND2X1 AND_tmp184 (.Y(ttmp184),.A(N1280),.B(N3018));
AND2X1 AND_tmp185 (.Y(N3505),.A(N468),.B(ttmp184));
AND2X1 AND_tmp186 (.Y(ttmp186),.A(N1280),.B(N3020));
AND2X1 AND_tmp187 (.Y(N3506),.A(N422),.B(ttmp186));
AND2X1 AND_tmp188 (.Y(ttmp188),.A(N1280),.B(N3022));
AND2X1 AND_tmp189 (.Y(N3507),.A(N435),.B(ttmp188));
AND2X1 AND2_551 (.Y(N3508),.A(N1685),.B(N3015));
AND2X1 AND2_552 (.Y(N3509),.A(N1685),.B(N3017));
AND2X1 AND2_553 (.Y(N3510),.A(N1685),.B(N3019));
AND2X1 AND2_554 (.Y(N3511),.A(N1685),.B(N3021));
NAND2X1 NAND2_555 (.Y(N3512),.A(N1923),.B(N3031));
NAND2X1 NAND2_556 (.Y(N3513),.A(N1920),.B(N3032));
NAND2X1 NAND2_557 (.Y(N3514),.A(N1929),.B(N3033));
NAND2X1 NAND2_558 (.Y(N3515),.A(N1926),.B(N3034));
NAND2X1 NAND2_559 (.Y(N3558),.A(N1947),.B(N3141));
NAND2X1 NAND2_560 (.Y(N3559),.A(N1944),.B(N3142));
NAND2X1 NAND2_561 (.Y(N3560),.A(N1953),.B(N3143));
NAND2X1 NAND2_562 (.Y(N3561),.A(N1950),.B(N3144));
NAND2X1 NAND2_563 (.Y(N3562),.A(N1959),.B(N3145));
NAND2X1 NAND2_564 (.Y(N3563),.A(N1956),.B(N3146));
BUFX1 BUFF1_565 (.Y(N3604),.A(N3191));
NAND2X1 NAND2_566 (.Y(N3605),.A(N1935),.B(N3194));
NAND2X1 NAND2_567 (.Y(N3606),.A(N1932),.B(N3195));
NAND2X1 NAND2_568 (.Y(N3607),.A(N1941),.B(N3196));
NAND2X1 NAND2_569 (.Y(N3608),.A(N1938),.B(N3197));
NAND2X1 NAND2_570 (.Y(N3609),.A(N1965),.B(N3198));
NAND2X1 NAND2_571 (.Y(N3610),.A(N1962),.B(N3199));
INVX1 NOT1_572 (.Y(N3613),.A(N3191));
AND2X1 AND2_573 (.Y(N3614),.A(N2882),.B(N2891));
AND2X1 AND2_574 (.Y(N3615),.A(N1482),.B(N2891));
AND2X1 AND_tmp190 (.Y(ttmp190),.A(N2653),.B(N1173));
AND2X1 AND_tmp191 (.Y(N3616),.A(N200),.B(ttmp190));
AND2X1 AND_tmp192 (.Y(ttmp192),.A(N2653),.B(N1173));
AND2X1 AND_tmp193 (.Y(N3617),.A(N203),.B(ttmp192));
AND2X1 AND_tmp194 (.Y(ttmp194),.A(N2653),.B(N1173));
AND2X1 AND_tmp195 (.Y(N3618),.A(N197),.B(ttmp194));
AND2X1 AND_tmp196 (.Y(ttmp196),.A(N2653),.B(N1173));
AND2X1 AND_tmp197 (.Y(N3619),.A(N194),.B(ttmp196));
AND2X1 AND_tmp198 (.Y(ttmp198),.A(N2653),.B(N1173));
AND2X1 AND_tmp199 (.Y(N3620),.A(N191),.B(ttmp198));
AND2X1 AND_tmp200 (.Y(ttmp200),.A(N2681),.B(N1197));
AND2X1 AND_tmp201 (.Y(N3621),.A(N182),.B(ttmp200));
AND2X1 AND_tmp202 (.Y(ttmp202),.A(N2681),.B(N1197));
AND2X1 AND_tmp203 (.Y(N3622),.A(N188),.B(ttmp202));
AND2X1 AND_tmp204 (.Y(ttmp204),.A(N2681),.B(N1197));
AND2X1 AND_tmp205 (.Y(N3623),.A(N155),.B(ttmp204));
AND2X1 AND_tmp206 (.Y(ttmp206),.A(N2681),.B(N1197));
AND2X1 AND_tmp207 (.Y(N3624),.A(N149),.B(ttmp206));
AND2X1 AND2_584 (.Y(N3625),.A(N2882),.B(N2891));
AND2X1 AND2_585 (.Y(N3626),.A(N1482),.B(N2891));
AND2X1 AND_tmp208 (.Y(ttmp208),.A(N2728),.B(N1235));
AND2X1 AND_tmp209 (.Y(N3627),.A(N200),.B(ttmp208));
AND2X1 AND_tmp210 (.Y(ttmp210),.A(N2728),.B(N1235));
AND2X1 AND_tmp211 (.Y(N3628),.A(N203),.B(ttmp210));
AND2X1 AND_tmp212 (.Y(ttmp212),.A(N2728),.B(N1235));
AND2X1 AND_tmp213 (.Y(N3629),.A(N197),.B(ttmp212));
AND2X1 AND_tmp214 (.Y(ttmp214),.A(N2728),.B(N1235));
AND2X1 AND_tmp215 (.Y(N3630),.A(N194),.B(ttmp214));
AND2X1 AND_tmp216 (.Y(ttmp216),.A(N2728),.B(N1235));
AND2X1 AND_tmp217 (.Y(N3631),.A(N191),.B(ttmp216));
AND2X1 AND_tmp218 (.Y(ttmp218),.A(N2756),.B(N1259));
AND2X1 AND_tmp219 (.Y(N3632),.A(N182),.B(ttmp218));
AND2X1 AND_tmp220 (.Y(ttmp220),.A(N2756),.B(N1259));
AND2X1 AND_tmp221 (.Y(N3633),.A(N188),.B(ttmp220));
AND2X1 AND_tmp222 (.Y(ttmp222),.A(N2756),.B(N1259));
AND2X1 AND_tmp223 (.Y(N3634),.A(N155),.B(ttmp222));
AND2X1 AND_tmp224 (.Y(ttmp224),.A(N2756),.B(N1259));
AND2X1 AND_tmp225 (.Y(N3635),.A(N149),.B(ttmp224));
AND2X1 AND2_595 (.Y(N3636),.A(N2882),.B(N2891));
AND2X1 AND2_596 (.Y(N3637),.A(N1482),.B(N2891));
AND2X1 AND_tmp226 (.Y(ttmp226),.A(N3075),.B(N1743));
AND2X1 AND_tmp227 (.Y(N3638),.A(N109),.B(ttmp226));
AND2X1 AND2_598 (.Y(N3639),.A(N2882),.B(N2891));
AND2X1 AND2_599 (.Y(N3640),.A(N1482),.B(N2891));
AND2X1 AND_tmp228 (.Y(ttmp228),.A(N2779),.B(N1339));
AND2X1 AND_tmp229 (.Y(N3641),.A(N11),.B(ttmp228));
AND2X1 AND_tmp230 (.Y(ttmp230),.A(N3041),.B(N1709));
AND2X1 AND_tmp231 (.Y(N3642),.A(N109),.B(ttmp230));
AND2X1 AND_tmp232 (.Y(ttmp232),.A(N3041),.B(N1709));
AND2X1 AND_tmp233 (.Y(N3643),.A(N46),.B(ttmp232));
AND2X1 AND_tmp234 (.Y(ttmp234),.A(N3041),.B(N1709));
AND2X1 AND_tmp235 (.Y(N3644),.A(N100),.B(ttmp234));
AND2X1 AND_tmp236 (.Y(ttmp236),.A(N3041),.B(N1709));
AND2X1 AND_tmp237 (.Y(N3645),.A(N91),.B(ttmp236));
AND2X1 AND_tmp238 (.Y(ttmp238),.A(N3041),.B(N1709));
AND2X1 AND_tmp239 (.Y(N3646),.A(N43),.B(ttmp238));
AND2X1 AND_tmp240 (.Y(ttmp240),.A(N2779),.B(N1339));
AND2X1 AND_tmp241 (.Y(N3647),.A(N76),.B(ttmp240));
AND2X1 AND_tmp242 (.Y(ttmp242),.A(N2779),.B(N1339));
AND2X1 AND_tmp243 (.Y(N3648),.A(N73),.B(ttmp242));
AND2X1 AND_tmp244 (.Y(ttmp244),.A(N2779),.B(N1339));
AND2X1 AND_tmp245 (.Y(N3649),.A(N67),.B(ttmp244));
AND2X1 AND_tmp246 (.Y(ttmp246),.A(N2779),.B(N1339));
AND2X1 AND_tmp247 (.Y(N3650),.A(N14),.B(ttmp246));
AND2X1 AND_tmp248 (.Y(ttmp248),.A(N3075),.B(N1743));
AND2X1 AND_tmp249 (.Y(N3651),.A(N46),.B(ttmp248));
AND2X1 AND_tmp250 (.Y(ttmp250),.A(N3075),.B(N1743));
AND2X1 AND_tmp251 (.Y(N3652),.A(N100),.B(ttmp250));
AND2X1 AND_tmp252 (.Y(ttmp252),.A(N3075),.B(N1743));
AND2X1 AND_tmp253 (.Y(N3653),.A(N91),.B(ttmp252));
AND2X1 AND_tmp254 (.Y(ttmp254),.A(N3075),.B(N1743));
AND2X1 AND_tmp255 (.Y(N3654),.A(N43),.B(ttmp254));
AND2X1 AND_tmp256 (.Y(ttmp256),.A(N2801),.B(N1363));
AND2X1 AND_tmp257 (.Y(N3655),.A(N76),.B(ttmp256));
AND2X1 AND_tmp258 (.Y(ttmp258),.A(N2801),.B(N1363));
AND2X1 AND_tmp259 (.Y(N3656),.A(N73),.B(ttmp258));
AND2X1 AND_tmp260 (.Y(ttmp260),.A(N2801),.B(N1363));
AND2X1 AND_tmp261 (.Y(N3657),.A(N67),.B(ttmp260));
AND2X1 AND_tmp262 (.Y(ttmp262),.A(N2801),.B(N1363));
AND2X1 AND_tmp263 (.Y(N3658),.A(N14),.B(ttmp262));
AND2X1 AND_tmp264 (.Y(ttmp264),.A(N3119),.B(N1785));
AND2X1 AND_tmp265 (.Y(N3659),.A(N120),.B(ttmp264));
AND2X1 AND_tmp266 (.Y(ttmp266),.A(N2801),.B(N1363));
AND2X1 AND_tmp267 (.Y(N3660),.A(N11),.B(ttmp266));
AND2X1 AND_tmp268 (.Y(ttmp268),.A(N3097),.B(N1769));
AND2X1 AND_tmp269 (.Y(N3661),.A(N118),.B(ttmp268));
AND2X1 AND_tmp270 (.Y(ttmp270),.A(N2681),.B(N1197));
AND2X1 AND_tmp271 (.Y(N3662),.A(N176),.B(ttmp270));
AND2X1 AND_tmp272 (.Y(ttmp272),.A(N2756),.B(N1259));
AND2X1 AND_tmp273 (.Y(N3663),.A(N176),.B(ttmp272));
OR2X1 OR2_623 (.Y(N3664),.A(N2831),.B(N3401));
OR2X1 OR2_624 (.Y(N3665),.A(N2832),.B(N3402));
OR2X1 OR2_625 (.Y(N3666),.A(N2833),.B(N3403));
OR2X1 OR2_626 (.Y(N3667),.A(N2834),.B(N3404));
OR2X1 OR_tmp274 (.Y(ttmp274),.A(N3405),.B(N457));
OR2X1 OR_tmp275 (.Y(N3668),.A(N2835),.B(ttmp274));
OR2X1 OR_tmp276 (.Y(ttmp276),.A(N3406),.B(N468));
OR2X1 OR_tmp277 (.Y(N3669),.A(N2836),.B(ttmp276));
OR2X1 OR_tmp278 (.Y(ttmp278),.A(N3407),.B(N422));
OR2X1 OR_tmp279 (.Y(N3670),.A(N2837),.B(ttmp278));
OR2X1 OR_tmp280 (.Y(ttmp280),.A(N3408),.B(N435));
OR2X1 OR_tmp281 (.Y(N3671),.A(N2838),.B(ttmp280));
OR2X1 OR2_631 (.Y(N3672),.A(N2847),.B(N3409));
OR2X1 OR2_632 (.Y(N3673),.A(N2848),.B(N3410));
OR2X1 OR2_633 (.Y(N3674),.A(N2849),.B(N3411));
OR2X1 OR2_634 (.Y(N3675),.A(N2850),.B(N3412));
OR2X1 OR_tmp282 (.Y(ttmp282),.A(N3413),.B(N389));
OR2X1 OR_tmp283 (.Y(N3676),.A(N2851),.B(ttmp282));
OR2X1 OR_tmp284 (.Y(ttmp284),.A(N3414),.B(N400));
OR2X1 OR_tmp285 (.Y(N3677),.A(N2852),.B(ttmp284));
OR2X1 OR_tmp286 (.Y(ttmp286),.A(N3415),.B(N411));
OR2X1 OR_tmp287 (.Y(N3678),.A(N2853),.B(ttmp286));
OR2X1 OR_tmp288 (.Y(ttmp288),.A(N3416),.B(N374));
OR2X1 OR_tmp289 (.Y(N3679),.A(N2854),.B(ttmp288));
AND2X1 AND2_639 (.Y(N3680),.A(N289),.B(N2855));
AND2X1 AND2_640 (.Y(N3681),.A(N281),.B(N2855));
AND2X1 AND2_641 (.Y(N3682),.A(N273),.B(N2855));
AND2X1 AND2_642 (.Y(N3683),.A(N265),.B(N2855));
AND2X1 AND2_643 (.Y(N3684),.A(N257),.B(N2855));
AND2X1 AND2_644 (.Y(N3685),.A(N234),.B(N2861));
AND2X1 AND2_645 (.Y(N3686),.A(N226),.B(N2861));
AND2X1 AND2_646 (.Y(N3687),.A(N218),.B(N2861));
AND2X1 AND2_647 (.Y(N3688),.A(N210),.B(N2861));
AND2X1 AND2_648 (.Y(N3689),.A(N206),.B(N2861));
INVX1 NOT1_649 (.Y(N3691),.A(N2891));
OR2X1 OR2_650 (.Y(N3700),.A(N2907),.B(N3444));
OR2X1 OR2_651 (.Y(N3701),.A(N2908),.B(N3445));
OR2X1 OR2_652 (.Y(N3702),.A(N2909),.B(N3446));
OR2X1 OR_tmp290 (.Y(ttmp290),.A(N3448),.B(N479));
OR2X1 OR_tmp291 (.Y(N3703),.A(N2911),.B(ttmp290));
OR2X1 OR_tmp292 (.Y(ttmp292),.A(N3449),.B(N490));
OR2X1 OR_tmp293 (.Y(N3704),.A(N2912),.B(ttmp292));
OR2X1 OR2_655 (.Y(N3705),.A(N2910),.B(N3447));
OR2X1 OR2_656 (.Y(N3708),.A(N2919),.B(N3450));
OR2X1 OR2_657 (.Y(N3709),.A(N2921),.B(N3451));
OR2X1 OR2_658 (.Y(N3710),.A(N2922),.B(N3452));
OR2X1 OR_tmp294 (.Y(ttmp294),.A(N3453),.B(N503));
OR2X1 OR_tmp295 (.Y(N3711),.A(N2923),.B(ttmp294));
OR2X1 OR_tmp296 (.Y(ttmp296),.A(N3454),.B(N523));
OR2X1 OR_tmp297 (.Y(N3712),.A(N2924),.B(ttmp296));
OR2X1 OR_tmp298 (.Y(ttmp298),.A(N3455),.B(N534));
OR2X1 OR_tmp299 (.Y(N3713),.A(N2925),.B(ttmp298));
OR2X1 OR2_662 (.Y(N3715),.A(N2934),.B(N3459));
OR2X1 OR2_663 (.Y(N3716),.A(N2935),.B(N3460));
OR2X1 OR2_664 (.Y(N3717),.A(N2936),.B(N3461));
OR2X1 OR2_665 (.Y(N3718),.A(N2937),.B(N3462));
OR2X1 OR_tmp300 (.Y(ttmp300),.A(N3463),.B(N389));
OR2X1 OR_tmp301 (.Y(N3719),.A(N2938),.B(ttmp300));
OR2X1 OR_tmp302 (.Y(ttmp302),.A(N3464),.B(N400));
OR2X1 OR_tmp303 (.Y(N3720),.A(N2939),.B(ttmp302));
OR2X1 OR_tmp304 (.Y(ttmp304),.A(N3465),.B(N411));
OR2X1 OR_tmp305 (.Y(N3721),.A(N2940),.B(ttmp304));
OR2X1 OR_tmp306 (.Y(ttmp306),.A(N3466),.B(N374));
OR2X1 OR_tmp307 (.Y(N3722),.A(N2941),.B(ttmp306));
AND2X1 AND2_670 (.Y(N3723),.A(N369),.B(N2942));
AND2X1 AND2_671 (.Y(N3724),.A(N361),.B(N2942));
AND2X1 AND2_672 (.Y(N3725),.A(N351),.B(N2942));
AND2X1 AND2_673 (.Y(N3726),.A(N341),.B(N2942));
AND2X1 AND2_674 (.Y(N3727),.A(N324),.B(N2948));
AND2X1 AND2_675 (.Y(N3728),.A(N316),.B(N2948));
AND2X1 AND2_676 (.Y(N3729),.A(N308),.B(N2948));
AND2X1 AND2_677 (.Y(N3730),.A(N302),.B(N2948));
AND2X1 AND2_678 (.Y(N3731),.A(N293),.B(N2948));
OR2X1 OR2_679 (.Y(N3732),.A(N2942),.B(N2958));
AND2X1 AND2_680 (.Y(N3738),.A(N83),.B(N2964));
AND2X1 AND2_681 (.Y(N3739),.A(N87),.B(N2964));
AND2X1 AND2_682 (.Y(N3740),.A(N34),.B(N2964));
AND2X1 AND2_683 (.Y(N3741),.A(N34),.B(N2964));
OR2X1 OR2_684 (.Y(N3742),.A(N2979),.B(N3481));
OR2X1 OR2_685 (.Y(N3743),.A(N2981),.B(N3483));
OR2X1 OR2_686 (.Y(N3744),.A(N2982),.B(N3484));
OR2X1 OR_tmp308 (.Y(ttmp308),.A(N3485),.B(N503));
OR2X1 OR_tmp309 (.Y(N3745),.A(N2983),.B(ttmp308));
OR2X1 OR_tmp310 (.Y(ttmp310),.A(N3486),.B(N523));
OR2X1 OR_tmp311 (.Y(N3746),.A(N2985),.B(ttmp310));
OR2X1 OR_tmp312 (.Y(ttmp312),.A(N3487),.B(N534));
OR2X1 OR_tmp313 (.Y(N3747),.A(N2986),.B(ttmp312));
OR2X1 OR2_690 (.Y(N3748),.A(N2993),.B(N3488));
OR2X1 OR2_691 (.Y(N3749),.A(N2994),.B(N3489));
OR2X1 OR2_692 (.Y(N3750),.A(N2995),.B(N3490));
OR2X1 OR_tmp314 (.Y(ttmp314),.A(N3492),.B(N479));
OR2X1 OR_tmp315 (.Y(N3751),.A(N2997),.B(ttmp314));
OR2X1 OR_tmp316 (.Y(ttmp316),.A(N3493),.B(N490));
OR2X1 OR_tmp317 (.Y(N3752),.A(N2998),.B(ttmp316));
INVX1 NOT1_695 (.Y(N3753),.A(N3000));
INVX1 NOT1_696 (.Y(N3754),.A(N3003));
INVX1 NOT1_697 (.Y(N3755),.A(N3007));
INVX1 NOT1_698 (.Y(N3756),.A(N3010));
OR2X1 OR2_699 (.Y(N3757),.A(N3013),.B(N3502));
AND2X1 AND_tmp318 (.Y(ttmp318),.A(N446),.B(N3003));
AND2X1 AND_tmp319 (.Y(N3758),.A(N1315),.B(ttmp318));
OR2X1 OR2_701 (.Y(N3759),.A(N3014),.B(N3503));
AND2X1 AND_tmp320 (.Y(ttmp320),.A(N446),.B(N3010));
AND2X1 AND_tmp321 (.Y(N3760),.A(N1315),.B(ttmp320));
AND2X1 AND2_703 (.Y(N3761),.A(N1675),.B(N3000));
AND2X1 AND2_704 (.Y(N3762),.A(N1675),.B(N3007));
OR2X1 OR2_705 (.Y(N3763),.A(N3023),.B(N3504));
OR2X1 OR2_706 (.Y(N3764),.A(N3024),.B(N3505));
OR2X1 OR2_707 (.Y(N3765),.A(N3025),.B(N3506));
OR2X1 OR2_708 (.Y(N3766),.A(N3026),.B(N3507));
OR2X1 OR_tmp322 (.Y(ttmp322),.A(N3508),.B(N457));
OR2X1 OR_tmp323 (.Y(N3767),.A(N3027),.B(ttmp322));
OR2X1 OR_tmp324 (.Y(ttmp324),.A(N3509),.B(N468));
OR2X1 OR_tmp325 (.Y(N3768),.A(N3028),.B(ttmp324));
OR2X1 OR_tmp326 (.Y(ttmp326),.A(N3510),.B(N422));
OR2X1 OR_tmp327 (.Y(N3769),.A(N3029),.B(ttmp326));
OR2X1 OR_tmp328 (.Y(ttmp328),.A(N3511),.B(N435));
OR2X1 OR_tmp329 (.Y(N3770),.A(N3030),.B(ttmp328));
NAND2X1 NAND2_713 (.Y(N3771),.A(N3512),.B(N3513));
NAND2X1 NAND2_714 (.Y(N3775),.A(N3514),.B(N3515));
INVX1 NOT1_715 (.Y(N3779),.A(N3035));
INVX1 NOT1_716 (.Y(N3780),.A(N3038));
AND2X1 AND_tmp330 (.Y(ttmp330),.A(N3097),.B(N1769));
AND2X1 AND_tmp331 (.Y(N3781),.A(N117),.B(ttmp330));
AND2X1 AND_tmp332 (.Y(ttmp332),.A(N3097),.B(N1769));
AND2X1 AND_tmp333 (.Y(N3782),.A(N126),.B(ttmp332));
AND2X1 AND_tmp334 (.Y(ttmp334),.A(N3097),.B(N1769));
AND2X1 AND_tmp335 (.Y(N3783),.A(N127),.B(ttmp334));
AND2X1 AND_tmp336 (.Y(ttmp336),.A(N3097),.B(N1769));
AND2X1 AND_tmp337 (.Y(N3784),.A(N128),.B(ttmp336));
AND2X1 AND_tmp338 (.Y(ttmp338),.A(N3119),.B(N1785));
AND2X1 AND_tmp339 (.Y(N3785),.A(N131),.B(ttmp338));
AND2X1 AND_tmp340 (.Y(ttmp340),.A(N3119),.B(N1785));
AND2X1 AND_tmp341 (.Y(N3786),.A(N129),.B(ttmp340));
AND2X1 AND_tmp342 (.Y(ttmp342),.A(N3119),.B(N1785));
AND2X1 AND_tmp343 (.Y(N3787),.A(N119),.B(ttmp342));
AND2X1 AND_tmp344 (.Y(ttmp344),.A(N3119),.B(N1785));
AND2X1 AND_tmp345 (.Y(N3788),.A(N130),.B(ttmp344));
NAND2X1 NAND2_725 (.Y(N3789),.A(N3558),.B(N3559));
NAND2X1 NAND2_726 (.Y(N3793),.A(N3560),.B(N3561));
NAND2X1 NAND2_727 (.Y(N3797),.A(N3562),.B(N3563));
AND2X1 AND_tmp346 (.Y(ttmp346),.A(N3147),.B(N1800));
AND2X1 AND_tmp347 (.Y(N3800),.A(N122),.B(ttmp346));
AND2X1 AND_tmp348 (.Y(ttmp348),.A(N3147),.B(N1800));
AND2X1 AND_tmp349 (.Y(N3801),.A(N113),.B(ttmp348));
AND2X1 AND_tmp350 (.Y(ttmp350),.A(N3147),.B(N1800));
AND2X1 AND_tmp351 (.Y(N3802),.A(N53),.B(ttmp350));
AND2X1 AND_tmp352 (.Y(ttmp352),.A(N3147),.B(N1800));
AND2X1 AND_tmp353 (.Y(N3803),.A(N114),.B(ttmp352));
AND2X1 AND_tmp354 (.Y(ttmp354),.A(N3147),.B(N1800));
AND2X1 AND_tmp355 (.Y(N3804),.A(N115),.B(ttmp354));
AND2X1 AND_tmp356 (.Y(ttmp356),.A(N3169),.B(N1814));
AND2X1 AND_tmp357 (.Y(N3805),.A(N52),.B(ttmp356));
AND2X1 AND_tmp358 (.Y(ttmp358),.A(N3169),.B(N1814));
AND2X1 AND_tmp359 (.Y(N3806),.A(N112),.B(ttmp358));
AND2X1 AND_tmp360 (.Y(ttmp360),.A(N3169),.B(N1814));
AND2X1 AND_tmp361 (.Y(N3807),.A(N116),.B(ttmp360));
AND2X1 AND_tmp362 (.Y(ttmp362),.A(N3169),.B(N1814));
AND2X1 AND_tmp363 (.Y(N3808),.A(N121),.B(ttmp362));
AND2X1 AND_tmp364 (.Y(ttmp364),.A(N3169),.B(N1814));
AND2X1 AND_tmp365 (.Y(N3809),.A(N123),.B(ttmp364));
NAND2X1 NAND2_738 (.Y(N3810),.A(N3607),.B(N3608));
NAND2X1 NAND2_739 (.Y(N3813),.A(N3605),.B(N3606));
AND2X1 AND2_740 (.Y(N3816),.A(N3482),.B(N2984));
OR2X1 OR2_741 (.Y(N3819),.A(N2996),.B(N3491));
INVX1 NOT1_742 (.Y(N3822),.A(N3200));
NAND2X1 NAND2_743 (.Y(N3823),.A(N3200),.B(N3203));
NAND2X1 NAND2_744 (.Y(N3824),.A(N3609),.B(N3610));
INVX1 NOT1_745 (.Y(N3827),.A(N3456));
OR2X1 OR2_746 (.Y(N3828),.A(N3739),.B(N2970));
OR2X1 OR2_747 (.Y(N3829),.A(N3740),.B(N2971));
OR2X1 OR2_748 (.Y(N3830),.A(N3741),.B(N2972));
OR2X1 OR2_749 (.Y(N3831),.A(N3738),.B(N2969));
INVX1 NOT1_750 (.Y(N3834),.A(N3664));
INVX1 NOT1_751 (.Y(N3835),.A(N3665));
INVX1 NOT1_752 (.Y(N3836),.A(N3666));
INVX1 NOT1_753 (.Y(N3837),.A(N3667));
INVX1 NOT1_754 (.Y(N3838),.A(N3672));
INVX1 NOT1_755 (.Y(N3839),.A(N3673));
INVX1 NOT1_756 (.Y(N3840),.A(N3674));
INVX1 NOT1_757 (.Y(N3841),.A(N3675));
OR2X1 OR2_758 (.Y(N3842),.A(N3681),.B(N2868));
OR2X1 OR2_759 (.Y(N3849),.A(N3682),.B(N2869));
OR2X1 OR2_760 (.Y(N3855),.A(N3683),.B(N2870));
OR2X1 OR2_761 (.Y(N3861),.A(N3684),.B(N2871));
OR2X1 OR2_762 (.Y(N3867),.A(N3685),.B(N2872));
OR2X1 OR2_763 (.Y(N3873),.A(N3686),.B(N2873));
OR2X1 OR2_764 (.Y(N3881),.A(N3687),.B(N2874));
OR2X1 OR2_765 (.Y(N3887),.A(N3688),.B(N2875));
OR2X1 OR2_766 (.Y(N3893),.A(N3689),.B(N2876));
INVX1 NOT1_767 (.Y(N3908),.A(N3701));
INVX1 NOT1_768 (.Y(N3909),.A(N3702));
INVX1 NOT1_769 (.Y(N3911),.A(N3700));
INVX1 NOT1_770 (.Y(N3914),.A(N3708));
INVX1 NOT1_771 (.Y(N3915),.A(N3709));
INVX1 NOT1_772 (.Y(N3916),.A(N3710));
INVX1 NOT1_773 (.Y(N3917),.A(N3715));
INVX1 NOT1_774 (.Y(N3918),.A(N3716));
INVX1 NOT1_775 (.Y(N3919),.A(N3717));
INVX1 NOT1_776 (.Y(N3920),.A(N3718));
OR2X1 OR2_777 (.Y(N3921),.A(N3724),.B(N2955));
OR2X1 OR2_778 (.Y(N3927),.A(N3725),.B(N2956));
OR2X1 OR2_779 (.Y(N3933),.A(N3726),.B(N2957));
OR2X1 OR2_780 (.Y(N3942),.A(N3727),.B(N2959));
OR2X1 OR2_781 (.Y(N3948),.A(N3728),.B(N2960));
OR2X1 OR2_782 (.Y(N3956),.A(N3729),.B(N2961));
OR2X1 OR2_783 (.Y(N3962),.A(N3730),.B(N2962));
OR2X1 OR2_784 (.Y(N3968),.A(N3731),.B(N2963));
INVX1 NOT1_785 (.Y(N3975),.A(N3742));
INVX1 NOT1_786 (.Y(N3976),.A(N3743));
INVX1 NOT1_787 (.Y(N3977),.A(N3744));
INVX1 NOT1_788 (.Y(N3978),.A(N3749));
INVX1 NOT1_789 (.Y(N3979),.A(N3750));
AND2X1 AND_tmp366 (.Y(ttmp366),.A(N1292),.B(N3754));
AND2X1 AND_tmp367 (.Y(N3980),.A(N446),.B(ttmp366));
AND2X1 AND_tmp368 (.Y(ttmp368),.A(N1292),.B(N3756));
AND2X1 AND_tmp369 (.Y(N3981),.A(N446),.B(ttmp368));
AND2X1 AND2_792 (.Y(N3982),.A(N1271),.B(N3753));
AND2X1 AND2_793 (.Y(N3983),.A(N1271),.B(N3755));
INVX1 NOT1_794 (.Y(N3984),.A(N3757));
INVX1 NOT1_795 (.Y(N3987),.A(N3759));
INVX1 NOT1_796 (.Y(N3988),.A(N3763));
INVX1 NOT1_797 (.Y(N3989),.A(N3764));
INVX1 NOT1_798 (.Y(N3990),.A(N3765));
INVX1 NOT1_799 (.Y(N3991),.A(N3766));
AND2X1 AND_tmp370 (.Y(ttmp370),.A(N3119),.B(N3130));
AND2X1 AND_tmp371 (.Y(N3998),.A(N3456),.B(ttmp370));
OR2X1 OR2_801 (.Y(N4008),.A(N3723),.B(N2954));
OR2X1 OR2_802 (.Y(N4011),.A(N3680),.B(N2867));
INVX1 NOT1_803 (.Y(N4021),.A(N3748));
NAND2X1 NAND2_804 (.Y(N4024),.A(N1968),.B(N3822));
INVX1 NOT1_805 (.Y(N4027),.A(N3705));
AND2X1 AND2_806 (.Y(N4031),.A(N3828),.B(N1583));
AND2X1 AND_tmp372 (.Y(ttmp372),.A(N2882),.B(N3691));
AND2X1 AND_tmp373 (.Y(N4032),.A(N24),.B(ttmp372));
AND2X1 AND_tmp374 (.Y(ttmp374),.A(N1482),.B(N3691));
AND2X1 AND_tmp375 (.Y(N4033),.A(N25),.B(ttmp374));
AND2X1 AND_tmp376 (.Y(ttmp376),.A(N2882),.B(N3691));
AND2X1 AND_tmp377 (.Y(N4034),.A(N26),.B(ttmp376));
AND2X1 AND_tmp378 (.Y(ttmp378),.A(N1482),.B(N3691));
AND2X1 AND_tmp379 (.Y(N4035),.A(N81),.B(ttmp378));
AND2X1 AND2_811 (.Y(N4036),.A(N3829),.B(N1583));
AND2X1 AND_tmp380 (.Y(ttmp380),.A(N2882),.B(N3691));
AND2X1 AND_tmp381 (.Y(N4037),.A(N79),.B(ttmp380));
AND2X1 AND_tmp382 (.Y(ttmp382),.A(N1482),.B(N3691));
AND2X1 AND_tmp383 (.Y(N4038),.A(N23),.B(ttmp382));
AND2X1 AND_tmp384 (.Y(ttmp384),.A(N2882),.B(N3691));
AND2X1 AND_tmp385 (.Y(N4039),.A(N82),.B(ttmp384));
AND2X1 AND_tmp386 (.Y(ttmp386),.A(N1482),.B(N3691));
AND2X1 AND_tmp387 (.Y(N4040),.A(N80),.B(ttmp386));
AND2X1 AND2_816 (.Y(N4041),.A(N3830),.B(N1583));
AND2X1 AND2_817 (.Y(N4042),.A(N3831),.B(N1583));
AND2X1 AND2_818 (.Y(N4067),.A(N3732),.B(N514));
AND2X1 AND2_819 (.Y(N4080),.A(N514),.B(N3732));
AND2X1 AND2_820 (.Y(N4088),.A(N3834),.B(N3668));
AND2X1 AND2_821 (.Y(N4091),.A(N3835),.B(N3669));
AND2X1 AND2_822 (.Y(N4094),.A(N3836),.B(N3670));
AND2X1 AND2_823 (.Y(N4097),.A(N3837),.B(N3671));
AND2X1 AND2_824 (.Y(N4100),.A(N3838),.B(N3676));
AND2X1 AND2_825 (.Y(N4103),.A(N3839),.B(N3677));
AND2X1 AND2_826 (.Y(N4106),.A(N3840),.B(N3678));
AND2X1 AND2_827 (.Y(N4109),.A(N3841),.B(N3679));
AND2X1 AND2_828 (.Y(N4144),.A(N3908),.B(N3703));
AND2X1 AND2_829 (.Y(N4147),.A(N3909),.B(N3704));
BUFX1 BUFF1_830 (.Y(N4150),.A(N3705));
AND2X1 AND2_831 (.Y(N4153),.A(N3914),.B(N3711));
AND2X1 AND2_832 (.Y(N4156),.A(N3915),.B(N3712));
AND2X1 AND2_833 (.Y(N4159),.A(N3916),.B(N3713));
OR2X1 OR2_834 (.Y(N4183),.A(N3758),.B(N3980));
OR2X1 OR2_835 (.Y(N4184),.A(N3760),.B(N3981));
OR2X1 OR_tmp388 (.Y(ttmp388),.A(N3982),.B(N446));
OR2X1 OR_tmp389 (.Y(N4185),.A(N3761),.B(ttmp388));
OR2X1 OR_tmp390 (.Y(ttmp390),.A(N3983),.B(N446));
OR2X1 OR_tmp391 (.Y(N4186),.A(N3762),.B(ttmp390));
INVX1 NOT1_838 (.Y(N4188),.A(N3771));
INVX1 NOT1_839 (.Y(N4191),.A(N3775));
AND2X1 AND_tmp392 (.Y(ttmp392),.A(N3771),.B(N3035));
AND2X1 AND_tmp393 (.Y(N4196),.A(N3775),.B(ttmp392));
AND2X1 AND_tmp394 (.Y(ttmp394),.A(N3119),.B(N3130));
AND2X1 AND_tmp395 (.Y(N4197),.A(N3987),.B(ttmp394));
AND2X1 AND2_842 (.Y(N4198),.A(N3920),.B(N3722));
INVX1 NOT1_843 (.Y(N4199),.A(N3816));
INVX1 NOT1_844 (.Y(N4200),.A(N3789));
INVX1 NOT1_845 (.Y(N4203),.A(N3793));
BUFX1 BUFF1_846 (.Y(N4206),.A(N3797));
BUFX1 BUFF1_847 (.Y(N4209),.A(N3797));
BUFX1 BUFF1_848 (.Y(N4212),.A(N3732));
BUFX1 BUFF1_849 (.Y(N4215),.A(N3732));
BUFX1 BUFF1_850 (.Y(N4219),.A(N3732));
INVX1 NOT1_851 (.Y(N4223),.A(N3810));
INVX1 NOT1_852 (.Y(N4224),.A(N3813));
AND2X1 AND2_853 (.Y(N4225),.A(N3918),.B(N3720));
AND2X1 AND2_854 (.Y(N4228),.A(N3919),.B(N3721));
AND2X1 AND2_855 (.Y(N4231),.A(N3991),.B(N3770));
AND2X1 AND2_856 (.Y(N4234),.A(N3917),.B(N3719));
AND2X1 AND2_857 (.Y(N4237),.A(N3989),.B(N3768));
AND2X1 AND2_858 (.Y(N4240),.A(N3990),.B(N3769));
AND2X1 AND2_859 (.Y(N4243),.A(N3988),.B(N3767));
AND2X1 AND2_860 (.Y(N4246),.A(N3976),.B(N3746));
AND2X1 AND2_861 (.Y(N4249),.A(N3977),.B(N3747));
AND2X1 AND2_862 (.Y(N4252),.A(N3975),.B(N3745));
AND2X1 AND2_863 (.Y(N4255),.A(N3978),.B(N3751));
AND2X1 AND2_864 (.Y(N4258),.A(N3979),.B(N3752));
INVX1 NOT1_865 (.Y(N4263),.A(N3819));
NAND2X1 NAND2_866 (.Y(N4264),.A(N4024),.B(N3823));
INVX1 NOT1_867 (.Y(N4267),.A(N3824));
AND2X1 AND2_868 (.Y(N4268),.A(N446),.B(N3893));
INVX1 NOT1_869 (.Y(N4269),.A(N3911));
INVX1 NOT1_870 (.Y(N4270),.A(N3984));
AND2X1 AND2_871 (.Y(N4271),.A(N3893),.B(N446));
INVX1 NOT1_872 (.Y(N4272),.A(N4031));
OR2X1 OR_tmp396 (.Y(ttmp396),.A(N3614),.B(N3615));
OR2X1 OR_tmp397 (.Y(ttmp397),.A(N4032),.B(ttmp396));
OR2X1 OR_tmp398 (.Y(N4273),.A(N4033),.B(ttmp397));
OR2X1 OR_tmp399 (.Y(ttmp399),.A(N3625),.B(N3626));
OR2X1 OR_tmp400 (.Y(ttmp400),.A(N4034),.B(ttmp399));
OR2X1 OR_tmp401 (.Y(N4274),.A(N4035),.B(ttmp400));
INVX1 NOT1_875 (.Y(N4275),.A(N4036));
OR2X1 OR_tmp402 (.Y(ttmp402),.A(N3636),.B(N3637));
OR2X1 OR_tmp403 (.Y(ttmp403),.A(N4037),.B(ttmp402));
OR2X1 OR_tmp404 (.Y(N4276),.A(N4038),.B(ttmp403));
OR2X1 OR_tmp405 (.Y(ttmp405),.A(N3639),.B(N3640));
OR2X1 OR_tmp406 (.Y(ttmp406),.A(N4039),.B(ttmp405));
OR2X1 OR_tmp407 (.Y(N4277),.A(N4040),.B(ttmp406));
INVX1 NOT1_878 (.Y(N4278),.A(N4041));
INVX1 NOT1_879 (.Y(N4279),.A(N4042));
AND2X1 AND2_880 (.Y(N4280),.A(N3887),.B(N457));
AND2X1 AND2_881 (.Y(N4284),.A(N3881),.B(N468));
AND2X1 AND2_882 (.Y(N4290),.A(N422),.B(N3873));
AND2X1 AND2_883 (.Y(N4297),.A(N3867),.B(N435));
AND2X1 AND2_884 (.Y(N4298),.A(N3861),.B(N389));
AND2X1 AND2_885 (.Y(N4301),.A(N3855),.B(N400));
AND2X1 AND2_886 (.Y(N4305),.A(N3849),.B(N411));
AND2X1 AND2_887 (.Y(N4310),.A(N3842),.B(N374));
AND2X1 AND2_888 (.Y(N4316),.A(N457),.B(N3887));
AND2X1 AND2_889 (.Y(N4320),.A(N468),.B(N3881));
AND2X1 AND2_890 (.Y(N4325),.A(N422),.B(N3873));
AND2X1 AND2_891 (.Y(N4331),.A(N435),.B(N3867));
AND2X1 AND2_892 (.Y(N4332),.A(N389),.B(N3861));
AND2X1 AND2_893 (.Y(N4336),.A(N400),.B(N3855));
AND2X1 AND2_894 (.Y(N4342),.A(N411),.B(N3849));
AND2X1 AND2_895 (.Y(N4349),.A(N374),.B(N3842));
INVX1 NOT1_896 (.Y(N4357),.A(N3968));
INVX1 NOT1_897 (.Y(N4364),.A(N3962));
BUFX1 BUFF1_898 (.Y(N4375),.A(N3962));
AND2X1 AND2_899 (.Y(N4379),.A(N3956),.B(N479));
AND2X1 AND2_900 (.Y(N4385),.A(N490),.B(N3948));
AND2X1 AND2_901 (.Y(N4392),.A(N3942),.B(N503));
AND2X1 AND2_902 (.Y(N4396),.A(N3933),.B(N523));
AND2X1 AND2_903 (.Y(N4400),.A(N3927),.B(N534));
INVX1 NOT1_904 (.Y(N4405),.A(N3921));
BUFX1 BUFF1_905 (.Y(N4412),.A(N3921));
INVX1 NOT1_906 (.Y(N4418),.A(N3968));
INVX1 NOT1_907 (.Y(N4425),.A(N3962));
BUFX1 BUFF1_908 (.Y(N4436),.A(N3962));
AND2X1 AND2_909 (.Y(N4440),.A(N479),.B(N3956));
AND2X1 AND2_910 (.Y(N4445),.A(N490),.B(N3948));
AND2X1 AND2_911 (.Y(N4451),.A(N503),.B(N3942));
AND2X1 AND2_912 (.Y(N4456),.A(N523),.B(N3933));
AND2X1 AND2_913 (.Y(N4462),.A(N534),.B(N3927));
BUFX1 BUFF1_914 (.Y(N4469),.A(N3921));
INVX1 NOT1_915 (.Y(N4477),.A(N3921));
BUFX1 BUFF1_916 (.Y(N4512),.A(N3968));
INVX1 NOT1_917 (.Y(N4515),.A(N4183));
INVX1 NOT1_918 (.Y(N4516),.A(N4184));
INVX1 NOT1_919 (.Y(N4521),.A(N4008));
INVX1 NOT1_920 (.Y(N4523),.A(N4011));
INVX1 NOT1_921 (.Y(N4524),.A(N4198));
INVX1 NOT1_922 (.Y(N4532),.A(N3984));
AND2X1 AND_tmp408 (.Y(ttmp408),.A(N3169),.B(N3180));
AND2X1 AND_tmp409 (.Y(N4547),.A(N3911),.B(ttmp408));
BUFX1 BUFF1_924 (.Y(N4548),.A(N3893));
BUFX1 BUFF1_925 (.Y(N4551),.A(N3887));
BUFX1 BUFF1_926 (.Y(N4554),.A(N3881));
BUFX1 BUFF1_927 (.Y(N4557),.A(N3873));
BUFX1 BUFF1_928 (.Y(N4560),.A(N3867));
BUFX1 BUFF1_929 (.Y(N4563),.A(N3861));
BUFX1 BUFF1_930 (.Y(N4566),.A(N3855));
BUFX1 BUFF1_931 (.Y(N4569),.A(N3849));
BUFX1 BUFF1_932 (.Y(N4572),.A(N3842));
NOR2X1 NOR2_933 (.Y(N4575),.A(N422),.B(N3873));
BUFX1 BUFF1_934 (.Y(N4578),.A(N3893));
BUFX1 BUFF1_935 (.Y(N4581),.A(N3887));
BUFX1 BUFF1_936 (.Y(N4584),.A(N3881));
BUFX1 BUFF1_937 (.Y(N4587),.A(N3867));
BUFX1 BUFF1_938 (.Y(N4590),.A(N3861));
BUFX1 BUFF1_939 (.Y(N4593),.A(N3855));
BUFX1 BUFF1_940 (.Y(N4596),.A(N3849));
BUFX1 BUFF1_941 (.Y(N4599),.A(N3873));
BUFX1 BUFF1_942 (.Y(N4602),.A(N3842));
NOR2X1 NOR2_943 (.Y(N4605),.A(N422),.B(N3873));
NOR2X1 NOR2_944 (.Y(N4608),.A(N374),.B(N3842));
BUFX1 BUFF1_945 (.Y(N4611),.A(N3956));
BUFX1 BUFF1_946 (.Y(N4614),.A(N3948));
BUFX1 BUFF1_947 (.Y(N4617),.A(N3942));
BUFX1 BUFF1_948 (.Y(N4621),.A(N3933));
BUFX1 BUFF1_949 (.Y(N4624),.A(N3927));
NOR2X1 NOR2_950 (.Y(N4627),.A(N490),.B(N3948));
BUFX1 BUFF1_951 (.Y(N4630),.A(N3956));
BUFX1 BUFF1_952 (.Y(N4633),.A(N3942));
BUFX1 BUFF1_953 (.Y(N4637),.A(N3933));
BUFX1 BUFF1_954 (.Y(N4640),.A(N3927));
BUFX1 BUFF1_955 (.Y(N4643),.A(N3948));
NOR2X1 NOR2_956 (.Y(N4646),.A(N490),.B(N3948));
BUFX1 BUFF1_957 (.Y(N4649),.A(N3927));
BUFX1 BUFF1_958 (.Y(N4652),.A(N3933));
BUFX1 BUFF1_959 (.Y(N4655),.A(N3921));
BUFX1 BUFF1_960 (.Y(N4658),.A(N3942));
BUFX1 BUFF1_961 (.Y(N4662),.A(N3956));
BUFX1 BUFF1_962 (.Y(N4665),.A(N3948));
BUFX1 BUFF1_963 (.Y(N4668),.A(N3968));
BUFX1 BUFF1_964 (.Y(N4671),.A(N3962));
BUFX1 BUFF1_965 (.Y(N4674),.A(N3873));
BUFX1 BUFF1_966 (.Y(N4677),.A(N3867));
BUFX1 BUFF1_967 (.Y(N4680),.A(N3887));
BUFX1 BUFF1_968 (.Y(N4683),.A(N3881));
BUFX1 BUFF1_969 (.Y(N4686),.A(N3893));
BUFX1 BUFF1_970 (.Y(N4689),.A(N3849));
BUFX1 BUFF1_971 (.Y(N4692),.A(N3842));
BUFX1 BUFF1_972 (.Y(N4695),.A(N3861));
BUFX1 BUFF1_973 (.Y(N4698),.A(N3855));
NAND2X1 NAND2_974 (.Y(N4701),.A(N3813),.B(N4223));
NAND2X1 NAND2_975 (.Y(N4702),.A(N3810),.B(N4224));
INVX1 NOT1_976 (.Y(N4720),.A(N4021));
NAND2X1 NAND2_977 (.Y(N4721),.A(N4021),.B(N4263));
INVX1 NOT1_978 (.Y(N4724),.A(N4147));
INVX1 NOT1_979 (.Y(N4725),.A(N4144));
INVX1 NOT1_980 (.Y(N4726),.A(N4159));
INVX1 NOT1_981 (.Y(N4727),.A(N4156));
INVX1 NOT1_982 (.Y(N4728),.A(N4153));
INVX1 NOT1_983 (.Y(N4729),.A(N4097));
INVX1 NOT1_984 (.Y(N4730),.A(N4094));
INVX1 NOT1_985 (.Y(N4731),.A(N4091));
INVX1 NOT1_986 (.Y(N4732),.A(N4088));
INVX1 NOT1_987 (.Y(N4733),.A(N4109));
INVX1 NOT1_988 (.Y(N4734),.A(N4106));
INVX1 NOT1_989 (.Y(N4735),.A(N4103));
INVX1 NOT1_990 (.Y(N4736),.A(N4100));
AND2X1 AND2_991 (.Y(N4737),.A(N4273),.B(N2877));
AND2X1 AND2_992 (.Y(N4738),.A(N4274),.B(N2877));
AND2X1 AND2_993 (.Y(N4739),.A(N4276),.B(N2877));
AND2X1 AND2_994 (.Y(N4740),.A(N4277),.B(N2877));
AND2X1 AND_tmp410 (.Y(ttmp410),.A(N1758),.B(N1755));
AND2X1 AND_tmp411 (.Y(N4741),.A(N4150),.B(ttmp410));
INVX1 NOT1_996 (.Y(N4855),.A(N4212));
NAND2X1 NAND2_997 (.Y(N4856),.A(N4212),.B(N2712));
NAND2X1 NAND2_998 (.Y(N4908),.A(N4215),.B(N2718));
INVX1 NOT1_999 (.Y(N4909),.A(N4215));
AND2X1 AND2_1000 (.Y(N4939),.A(N4515),.B(N4185));
AND2X1 AND2_1001 (.Y(N4942),.A(N4516),.B(N4186));
INVX1 NOT1_1002 (.Y(N4947),.A(N4219));
AND2X1 AND_tmp412 (.Y(ttmp412),.A(N3775),.B(N3779));
AND2X1 AND_tmp413 (.Y(N4953),.A(N4188),.B(ttmp412));
AND2X1 AND_tmp414 (.Y(ttmp414),.A(N4191),.B(N3780));
AND2X1 AND_tmp415 (.Y(N4954),.A(N3771),.B(ttmp414));
AND2X1 AND_tmp416 (.Y(ttmp416),.A(N4188),.B(N3038));
AND2X1 AND_tmp417 (.Y(N4955),.A(N4191),.B(ttmp416));
AND2X1 AND_tmp418 (.Y(ttmp418),.A(N3097),.B(N3108));
AND2X1 AND_tmp419 (.Y(N4956),.A(N4109),.B(ttmp418));
AND2X1 AND_tmp420 (.Y(ttmp420),.A(N3097),.B(N3108));
AND2X1 AND_tmp421 (.Y(N4957),.A(N4106),.B(ttmp420));
AND2X1 AND_tmp422 (.Y(ttmp422),.A(N3097),.B(N3108));
AND2X1 AND_tmp423 (.Y(N4958),.A(N4103),.B(ttmp422));
AND2X1 AND_tmp424 (.Y(ttmp424),.A(N3097),.B(N3108));
AND2X1 AND_tmp425 (.Y(N4959),.A(N4100),.B(ttmp424));
AND2X1 AND_tmp426 (.Y(ttmp426),.A(N3119),.B(N3130));
AND2X1 AND_tmp427 (.Y(N4960),.A(N4159),.B(ttmp426));
AND2X1 AND_tmp428 (.Y(ttmp428),.A(N3119),.B(N3130));
AND2X1 AND_tmp429 (.Y(N4961),.A(N4156),.B(ttmp428));
INVX1 NOT1_1012 (.Y(N4965),.A(N4225));
INVX1 NOT1_1013 (.Y(N4966),.A(N4228));
INVX1 NOT1_1014 (.Y(N4967),.A(N4231));
INVX1 NOT1_1015 (.Y(N4968),.A(N4234));
INVX1 NOT1_1016 (.Y(N4972),.A(N4246));
INVX1 NOT1_1017 (.Y(N4973),.A(N4249));
INVX1 NOT1_1018 (.Y(N4974),.A(N4252));
NAND2X1 NAND2_1019 (.Y(N4975),.A(N4252),.B(N4199));
INVX1 NOT1_1020 (.Y(N4976),.A(N4206));
INVX1 NOT1_1021 (.Y(N4977),.A(N4209));
AND2X1 AND_tmp430 (.Y(ttmp430),.A(N3789),.B(N4206));
AND2X1 AND_tmp431 (.Y(N4978),.A(N3793),.B(ttmp430));
AND2X1 AND_tmp432 (.Y(ttmp432),.A(N4200),.B(N4209));
AND2X1 AND_tmp433 (.Y(N4979),.A(N4203),.B(ttmp432));
AND2X1 AND_tmp434 (.Y(ttmp434),.A(N3147),.B(N3158));
AND2X1 AND_tmp435 (.Y(N4980),.A(N4097),.B(ttmp434));
AND2X1 AND_tmp436 (.Y(ttmp436),.A(N3147),.B(N3158));
AND2X1 AND_tmp437 (.Y(N4981),.A(N4094),.B(ttmp436));
AND2X1 AND_tmp438 (.Y(ttmp438),.A(N3147),.B(N3158));
AND2X1 AND_tmp439 (.Y(N4982),.A(N4091),.B(ttmp438));
AND2X1 AND_tmp440 (.Y(ttmp440),.A(N3147),.B(N3158));
AND2X1 AND_tmp441 (.Y(N4983),.A(N4088),.B(ttmp440));
AND2X1 AND_tmp442 (.Y(ttmp442),.A(N3169),.B(N3180));
AND2X1 AND_tmp443 (.Y(N4984),.A(N4153),.B(ttmp442));
AND2X1 AND_tmp444 (.Y(ttmp444),.A(N3169),.B(N3180));
AND2X1 AND_tmp445 (.Y(N4985),.A(N4147),.B(ttmp444));
AND2X1 AND_tmp446 (.Y(ttmp446),.A(N3169),.B(N3180));
AND2X1 AND_tmp447 (.Y(N4986),.A(N4144),.B(ttmp446));
AND2X1 AND_tmp448 (.Y(ttmp448),.A(N3169),.B(N3180));
AND2X1 AND_tmp449 (.Y(N4987),.A(N4150),.B(ttmp448));
NAND2X1 NAND2_1032 (.Y(N5049),.A(N4701),.B(N4702));
INVX1 NOT1_1033 (.Y(N5052),.A(N4237));
INVX1 NOT1_1034 (.Y(N5053),.A(N4240));
INVX1 NOT1_1035 (.Y(N5054),.A(N4243));
INVX1 NOT1_1036 (.Y(N5055),.A(N4255));
INVX1 NOT1_1037 (.Y(N5056),.A(N4258));
NAND2X1 NAND2_1038 (.Y(N5057),.A(N3819),.B(N4720));
INVX1 NOT1_1039 (.Y(N5058),.A(N4264));
NAND2X1 NAND2_1040 (.Y(N5059),.A(N4264),.B(N4267));
AND2X1 AND_tmp450 (.Y(ttmp450),.A(N4269),.B(N4027));
AND2X1 AND_tmp451 (.Y(ttmp451),.A(N4724),.B(ttmp450));
AND2X1 AND_tmp452 (.Y(N5060),.A(N4725),.B(ttmp451));
AND2X1 AND_tmp453 (.Y(ttmp453),.A(N3827),.B(N4728));
AND2X1 AND_tmp454 (.Y(ttmp454),.A(N4726),.B(ttmp453));
AND2X1 AND_tmp455 (.Y(N5061),.A(N4727),.B(ttmp454));
AND2X1 AND_tmp456 (.Y(ttmp456),.A(N4731),.B(N4732));
AND2X1 AND_tmp457 (.Y(ttmp457),.A(N4729),.B(ttmp456));
AND2X1 AND_tmp458 (.Y(N5062),.A(N4730),.B(ttmp457));
AND2X1 AND_tmp459 (.Y(ttmp459),.A(N4735),.B(N4736));
AND2X1 AND_tmp460 (.Y(ttmp460),.A(N4733),.B(ttmp459));
AND2X1 AND_tmp461 (.Y(N5063),.A(N4734),.B(ttmp460));
AND2X1 AND2_1045 (.Y(N5065),.A(N4357),.B(N4375));
AND2X1 AND_tmp462 (.Y(ttmp462),.A(N4357),.B(N4379));
AND2X1 AND_tmp463 (.Y(N5066),.A(N4364),.B(ttmp462));
AND2X1 AND2_1047 (.Y(N5067),.A(N4418),.B(N4436));
AND2X1 AND_tmp464 (.Y(ttmp464),.A(N4418),.B(N4440));
AND2X1 AND_tmp465 (.Y(N5068),.A(N4425),.B(ttmp464));
INVX1 NOT1_1049 (.Y(N5069),.A(N4548));
NAND2X1 NAND2_1050 (.Y(N5070),.A(N4548),.B(N2628));
INVX1 NOT1_1051 (.Y(N5071),.A(N4551));
NAND2X1 NAND2_1052 (.Y(N5072),.A(N4551),.B(N2629));
INVX1 NOT1_1053 (.Y(N5073),.A(N4554));
NAND2X1 NAND2_1054 (.Y(N5074),.A(N4554),.B(N2630));
INVX1 NOT1_1055 (.Y(N5075),.A(N4557));
NAND2X1 NAND2_1056 (.Y(N5076),.A(N4557),.B(N2631));
INVX1 NOT1_1057 (.Y(N5077),.A(N4560));
NAND2X1 NAND2_1058 (.Y(N5078),.A(N4560),.B(N2632));
INVX1 NOT1_1059 (.Y(N5079),.A(N4563));
NAND2X1 NAND2_1060 (.Y(N5080),.A(N4563),.B(N2633));
INVX1 NOT1_1061 (.Y(N5081),.A(N4566));
NAND2X1 NAND2_1062 (.Y(N5082),.A(N4566),.B(N2634));
INVX1 NOT1_1063 (.Y(N5083),.A(N4569));
NAND2X1 NAND2_1064 (.Y(N5084),.A(N4569),.B(N2635));
INVX1 NOT1_1065 (.Y(N5085),.A(N4572));
NAND2X1 NAND2_1066 (.Y(N5086),.A(N4572),.B(N2636));
INVX1 NOT1_1067 (.Y(N5087),.A(N4575));
NAND2X1 NAND2_1068 (.Y(N5088),.A(N4578),.B(N2638));
INVX1 NOT1_1069 (.Y(N5089),.A(N4578));
NAND2X1 NAND2_1070 (.Y(N5090),.A(N4581),.B(N2639));
INVX1 NOT1_1071 (.Y(N5091),.A(N4581));
NAND2X1 NAND2_1072 (.Y(N5092),.A(N4584),.B(N2640));
INVX1 NOT1_1073 (.Y(N5093),.A(N4584));
NAND2X1 NAND2_1074 (.Y(N5094),.A(N4587),.B(N2641));
INVX1 NOT1_1075 (.Y(N5095),.A(N4587));
NAND2X1 NAND2_1076 (.Y(N5096),.A(N4590),.B(N2642));
INVX1 NOT1_1077 (.Y(N5097),.A(N4590));
NAND2X1 NAND2_1078 (.Y(N5098),.A(N4593),.B(N2643));
INVX1 NOT1_1079 (.Y(N5099),.A(N4593));
NAND2X1 NAND2_1080 (.Y(N5100),.A(N4596),.B(N2644));
INVX1 NOT1_1081 (.Y(N5101),.A(N4596));
NAND2X1 NAND2_1082 (.Y(N5102),.A(N4599),.B(N2645));
INVX1 NOT1_1083 (.Y(N5103),.A(N4599));
NAND2X1 NAND2_1084 (.Y(N5104),.A(N4602),.B(N2646));
INVX1 NOT1_1085 (.Y(N5105),.A(N4602));
INVX1 NOT1_1086 (.Y(N5106),.A(N4611));
NAND2X1 NAND2_1087 (.Y(N5107),.A(N4611),.B(N2709));
INVX1 NOT1_1088 (.Y(N5108),.A(N4614));
NAND2X1 NAND2_1089 (.Y(N5109),.A(N4614),.B(N2710));
INVX1 NOT1_1090 (.Y(N5110),.A(N4617));
NAND2X1 NAND2_1091 (.Y(N5111),.A(N4617),.B(N2711));
NAND2X1 NAND2_1092 (.Y(N5112),.A(N1890),.B(N4855));
INVX1 NOT1_1093 (.Y(N5113),.A(N4621));
NAND2X1 NAND2_1094 (.Y(N5114),.A(N4621),.B(N2713));
INVX1 NOT1_1095 (.Y(N5115),.A(N4624));
NAND2X1 NAND2_1096 (.Y(N5116),.A(N4624),.B(N2714));
AND2X1 AND2_1097 (.Y(N5117),.A(N4364),.B(N4379));
AND2X1 AND2_1098 (.Y(N5118),.A(N4364),.B(N4379));
AND2X1 AND2_1099 (.Y(N5119),.A(N54),.B(N4405));
INVX1 NOT1_1100 (.Y(N5120),.A(N4627));
NAND2X1 NAND2_1101 (.Y(N5121),.A(N4630),.B(N2716));
INVX1 NOT1_1102 (.Y(N5122),.A(N4630));
NAND2X1 NAND2_1103 (.Y(N5123),.A(N4633),.B(N2717));
INVX1 NOT1_1104 (.Y(N5124),.A(N4633));
NAND2X1 NAND2_1105 (.Y(N5125),.A(N1908),.B(N4909));
NAND2X1 NAND2_1106 (.Y(N5126),.A(N4637),.B(N2719));
INVX1 NOT1_1107 (.Y(N5127),.A(N4637));
NAND2X1 NAND2_1108 (.Y(N5128),.A(N4640),.B(N2720));
INVX1 NOT1_1109 (.Y(N5129),.A(N4640));
NAND2X1 NAND2_1110 (.Y(N5130),.A(N4643),.B(N2721));
INVX1 NOT1_1111 (.Y(N5131),.A(N4643));
AND2X1 AND2_1112 (.Y(N5132),.A(N4425),.B(N4440));
AND2X1 AND2_1113 (.Y(N5133),.A(N4425),.B(N4440));
INVX1 NOT1_1114 (.Y(N5135),.A(N4649));
INVX1 NOT1_1115 (.Y(N5136),.A(N4652));
NAND2X1 NAND2_1116 (.Y(N5137),.A(N4655),.B(N4521));
INVX1 NOT1_1117 (.Y(N5138),.A(N4655));
INVX1 NOT1_1118 (.Y(N5139),.A(N4658));
NAND2X1 NAND2_1119 (.Y(N5140),.A(N4658),.B(N4947));
INVX1 NOT1_1120 (.Y(N5141),.A(N4674));
INVX1 NOT1_1121 (.Y(N5142),.A(N4677));
INVX1 NOT1_1122 (.Y(N5143),.A(N4680));
INVX1 NOT1_1123 (.Y(N5144),.A(N4683));
NAND2X1 NAND2_1124 (.Y(N5145),.A(N4686),.B(N4523));
INVX1 NOT1_1125 (.Y(N5146),.A(N4686));
NOR2X1 NOR2_1126 (.Y(N5147),.A(N4953),.B(N4196));
NOR2X1 NOR2_1127 (.Y(N5148),.A(N4954),.B(N4955));
INVX1 NOT1_1128 (.Y(N5150),.A(N4524));
NAND2X1 NAND2_1129 (.Y(N5153),.A(N4228),.B(N4965));
NAND2X1 NAND2_1130 (.Y(N5154),.A(N4225),.B(N4966));
NAND2X1 NAND2_1131 (.Y(N5155),.A(N4234),.B(N4967));
NAND2X1 NAND2_1132 (.Y(N5156),.A(N4231),.B(N4968));
INVX1 NOT1_1133 (.Y(N5157),.A(N4532));
NAND2X1 NAND2_1134 (.Y(N5160),.A(N4249),.B(N4972));
NAND2X1 NAND2_1135 (.Y(N5161),.A(N4246),.B(N4973));
NAND2X1 NAND2_1136 (.Y(N5162),.A(N3816),.B(N4974));
AND2X1 AND_tmp466 (.Y(ttmp466),.A(N3793),.B(N4976));
AND2X1 AND_tmp467 (.Y(N5163),.A(N4200),.B(ttmp466));
AND2X1 AND_tmp468 (.Y(ttmp468),.A(N4203),.B(N4977));
AND2X1 AND_tmp469 (.Y(N5164),.A(N3789),.B(ttmp468));
AND2X1 AND_tmp470 (.Y(ttmp470),.A(N3147),.B(N3158));
AND2X1 AND_tmp471 (.Y(N5165),.A(N4942),.B(ttmp470));
INVX1 NOT1_1140 (.Y(N5166),.A(N4512));
BUFX1 BUFF1_1141 (.Y(N5169),.A(N4290));
INVX1 NOT1_1142 (.Y(N5172),.A(N4605));
BUFX1 BUFF1_1143 (.Y(N5173),.A(N4325));
INVX1 NOT1_1144 (.Y(N5176),.A(N4608));
BUFX1 BUFF1_1145 (.Y(N5177),.A(N4349));
BUFX1 BUFF1_1146 (.Y(N5180),.A(N4405));
BUFX1 BUFF1_1147 (.Y(N5183),.A(N4357));
BUFX1 BUFF1_1148 (.Y(N5186),.A(N4357));
BUFX1 BUFF1_1149 (.Y(N5189),.A(N4364));
BUFX1 BUFF1_1150 (.Y(N5192),.A(N4364));
BUFX1 BUFF1_1151 (.Y(N5195),.A(N4385));
INVX1 NOT1_1152 (.Y(N5198),.A(N4646));
BUFX1 BUFF1_1153 (.Y(N5199),.A(N4418));
BUFX1 BUFF1_1154 (.Y(N5202),.A(N4425));
BUFX1 BUFF1_1155 (.Y(N5205),.A(N4445));
BUFX1 BUFF1_1156 (.Y(N5208),.A(N4418));
BUFX1 BUFF1_1157 (.Y(N5211),.A(N4425));
BUFX1 BUFF1_1158 (.Y(N5214),.A(N4477));
BUFX1 BUFF1_1159 (.Y(N5217),.A(N4469));
BUFX1 BUFF1_1160 (.Y(N5220),.A(N4477));
INVX1 NOT1_1161 (.Y(N5223),.A(N4662));
INVX1 NOT1_1162 (.Y(N5224),.A(N4665));
INVX1 NOT1_1163 (.Y(N5225),.A(N4668));
INVX1 NOT1_1164 (.Y(N5226),.A(N4671));
INVX1 NOT1_1165 (.Y(N5227),.A(N4689));
INVX1 NOT1_1166 (.Y(N5228),.A(N4692));
INVX1 NOT1_1167 (.Y(N5229),.A(N4695));
INVX1 NOT1_1168 (.Y(N5230),.A(N4698));
NAND2X1 NAND2_1169 (.Y(N5232),.A(N4240),.B(N5052));
NAND2X1 NAND2_1170 (.Y(N5233),.A(N4237),.B(N5053));
NAND2X1 NAND2_1171 (.Y(N5234),.A(N4258),.B(N5055));
NAND2X1 NAND2_1172 (.Y(N5235),.A(N4255),.B(N5056));
NAND2X1 NAND2_1173 (.Y(N5236),.A(N4721),.B(N5057));
NAND2X1 NAND2_1174 (.Y(N5239),.A(N3824),.B(N5058));
AND2X1 AND_tmp472 (.Y(ttmp472),.A(N5061),.B(N4270));
AND2X1 AND_tmp473 (.Y(N5240),.A(N5060),.B(ttmp472));
INVX1 NOT1_1176 (.Y(N5241),.A(N4939));
NAND2X1 NAND2_1177 (.Y(N5242),.A(N1824),.B(N5069));
NAND2X1 NAND2_1178 (.Y(N5243),.A(N1827),.B(N5071));
NAND2X1 NAND2_1179 (.Y(N5244),.A(N1830),.B(N5073));
NAND2X1 NAND2_1180 (.Y(N5245),.A(N1833),.B(N5075));
NAND2X1 NAND2_1181 (.Y(N5246),.A(N1836),.B(N5077));
NAND2X1 NAND2_1182 (.Y(N5247),.A(N1839),.B(N5079));
NAND2X1 NAND2_1183 (.Y(N5248),.A(N1842),.B(N5081));
NAND2X1 NAND2_1184 (.Y(N5249),.A(N1845),.B(N5083));
NAND2X1 NAND2_1185 (.Y(N5250),.A(N1848),.B(N5085));
NAND2X1 NAND2_1186 (.Y(N5252),.A(N1854),.B(N5089));
NAND2X1 NAND2_1187 (.Y(N5253),.A(N1857),.B(N5091));
NAND2X1 NAND2_1188 (.Y(N5254),.A(N1860),.B(N5093));
NAND2X1 NAND2_1189 (.Y(N5255),.A(N1863),.B(N5095));
NAND2X1 NAND2_1190 (.Y(N5256),.A(N1866),.B(N5097));
NAND2X1 NAND2_1191 (.Y(N5257),.A(N1869),.B(N5099));
NAND2X1 NAND2_1192 (.Y(N5258),.A(N1872),.B(N5101));
NAND2X1 NAND2_1193 (.Y(N5259),.A(N1875),.B(N5103));
NAND2X1 NAND2_1194 (.Y(N5260),.A(N1878),.B(N5105));
NAND2X1 NAND2_1195 (.Y(N5261),.A(N1881),.B(N5106));
NAND2X1 NAND2_1196 (.Y(N5262),.A(N1884),.B(N5108));
NAND2X1 NAND2_1197 (.Y(N5263),.A(N1887),.B(N5110));
NAND2X1 NAND2_1198 (.Y(N5264),.A(N5112),.B(N4856));
NAND2X1 NAND2_1199 (.Y(N5274),.A(N1893),.B(N5113));
NAND2X1 NAND2_1200 (.Y(N5275),.A(N1896),.B(N5115));
NAND2X1 NAND2_1201 (.Y(N5282),.A(N1902),.B(N5122));
NAND2X1 NAND2_1202 (.Y(N5283),.A(N1905),.B(N5124));
NAND2X1 NAND2_1203 (.Y(N5284),.A(N4908),.B(N5125));
NAND2X1 NAND2_1204 (.Y(N5298),.A(N1911),.B(N5127));
NAND2X1 NAND2_1205 (.Y(N5299),.A(N1914),.B(N5129));
NAND2X1 NAND2_1206 (.Y(N5300),.A(N1917),.B(N5131));
NAND2X1 NAND2_1207 (.Y(N5303),.A(N4652),.B(N5135));
NAND2X1 NAND2_1208 (.Y(N5304),.A(N4649),.B(N5136));
NAND2X1 NAND2_1209 (.Y(N5305),.A(N4008),.B(N5138));
NAND2X1 NAND2_1210 (.Y(N5306),.A(N4219),.B(N5139));
NAND2X1 NAND2_1211 (.Y(N5307),.A(N4677),.B(N5141));
NAND2X1 NAND2_1212 (.Y(N5308),.A(N4674),.B(N5142));
NAND2X1 NAND2_1213 (.Y(N5309),.A(N4683),.B(N5143));
NAND2X1 NAND2_1214 (.Y(N5310),.A(N4680),.B(N5144));
NAND2X1 NAND2_1215 (.Y(N5311),.A(N4011),.B(N5146));
INVX1 NOT1_1216 (.Y(N5312),.A(N5049));
NAND2X1 NAND2_1217 (.Y(N5315),.A(N5153),.B(N5154));
NAND2X1 NAND2_1218 (.Y(N5319),.A(N5155),.B(N5156));
NAND2X1 NAND2_1219 (.Y(N5324),.A(N5160),.B(N5161));
NAND2X1 NAND2_1220 (.Y(N5328),.A(N5162),.B(N4975));
NOR2X1 NOR2_1221 (.Y(N5331),.A(N5163),.B(N4978));
NOR2X1 NOR2_1222 (.Y(N5332),.A(N5164),.B(N4979));
OR2X1 OR2_1223 (.Y(N5346),.A(N4412),.B(N5119));
NAND2X1 NAND2_1224 (.Y(N5363),.A(N4665),.B(N5223));
NAND2X1 NAND2_1225 (.Y(N5364),.A(N4662),.B(N5224));
NAND2X1 NAND2_1226 (.Y(N5365),.A(N4671),.B(N5225));
NAND2X1 NAND2_1227 (.Y(N5366),.A(N4668),.B(N5226));
NAND2X1 NAND2_1228 (.Y(N5367),.A(N4692),.B(N5227));
NAND2X1 NAND2_1229 (.Y(N5368),.A(N4689),.B(N5228));
NAND2X1 NAND2_1230 (.Y(N5369),.A(N4698),.B(N5229));
NAND2X1 NAND2_1231 (.Y(N5370),.A(N4695),.B(N5230));
NAND2X1 NAND2_1232 (.Y(N5371),.A(N5148),.B(N5147));
BUFX1 BUFF1_1233 (.Y(N5374),.A(N4939));
NAND2X1 NAND2_1234 (.Y(N5377),.A(N5232),.B(N5233));
NAND2X1 NAND2_1235 (.Y(N5382),.A(N5234),.B(N5235));
NAND2X1 NAND2_1236 (.Y(N5385),.A(N5239),.B(N5059));
AND2X1 AND_tmp474 (.Y(ttmp474),.A(N5063),.B(N5241));
AND2X1 AND_tmp475 (.Y(N5388),.A(N5062),.B(ttmp474));
NAND2X1 NAND2_1238 (.Y(N5389),.A(N5242),.B(N5070));
NAND2X1 NAND2_1239 (.Y(N5396),.A(N5243),.B(N5072));
NAND2X1 NAND2_1240 (.Y(N5407),.A(N5244),.B(N5074));
NAND2X1 NAND2_1241 (.Y(N5418),.A(N5245),.B(N5076));
NAND2X1 NAND2_1242 (.Y(N5424),.A(N5246),.B(N5078));
NAND2X1 NAND2_1243 (.Y(N5431),.A(N5247),.B(N5080));
NAND2X1 NAND2_1244 (.Y(N5441),.A(N5248),.B(N5082));
NAND2X1 NAND2_1245 (.Y(N5452),.A(N5249),.B(N5084));
NAND2X1 NAND2_1246 (.Y(N5462),.A(N5250),.B(N5086));
INVX1 NOT1_1247 (.Y(N5469),.A(N5169));
NAND2X1 NAND2_1248 (.Y(N5470),.A(N5088),.B(N5252));
NAND2X1 NAND2_1249 (.Y(N5477),.A(N5090),.B(N5253));
NAND2X1 NAND2_1250 (.Y(N5488),.A(N5092),.B(N5254));
NAND2X1 NAND2_1251 (.Y(N5498),.A(N5094),.B(N5255));
NAND2X1 NAND2_1252 (.Y(N5506),.A(N5096),.B(N5256));
NAND2X1 NAND2_1253 (.Y(N5520),.A(N5098),.B(N5257));
NAND2X1 NAND2_1254 (.Y(N5536),.A(N5100),.B(N5258));
NAND2X1 NAND2_1255 (.Y(N5549),.A(N5102),.B(N5259));
NAND2X1 NAND2_1256 (.Y(N5555),.A(N5104),.B(N5260));
NAND2X1 NAND2_1257 (.Y(N5562),.A(N5261),.B(N5107));
NAND2X1 NAND2_1258 (.Y(N5573),.A(N5262),.B(N5109));
NAND2X1 NAND2_1259 (.Y(N5579),.A(N5263),.B(N5111));
NAND2X1 NAND2_1260 (.Y(N5595),.A(N5274),.B(N5114));
NAND2X1 NAND2_1261 (.Y(N5606),.A(N5275),.B(N5116));
NAND2X1 NAND2_1262 (.Y(N5616),.A(N5180),.B(N2715));
INVX1 NOT1_1263 (.Y(N5617),.A(N5180));
INVX1 NOT1_1264 (.Y(N5618),.A(N5183));
INVX1 NOT1_1265 (.Y(N5619),.A(N5186));
INVX1 NOT1_1266 (.Y(N5620),.A(N5189));
INVX1 NOT1_1267 (.Y(N5621),.A(N5192));
INVX1 NOT1_1268 (.Y(N5622),.A(N5195));
NAND2X1 NAND2_1269 (.Y(N5624),.A(N5121),.B(N5282));
NAND2X1 NAND2_1270 (.Y(N5634),.A(N5123),.B(N5283));
NAND2X1 NAND2_1271 (.Y(N5655),.A(N5126),.B(N5298));
NAND2X1 NAND2_1272 (.Y(N5671),.A(N5128),.B(N5299));
NAND2X1 NAND2_1273 (.Y(N5684),.A(N5130),.B(N5300));
INVX1 NOT1_1274 (.Y(N5690),.A(N5202));
INVX1 NOT1_1275 (.Y(N5691),.A(N5211));
NAND2X1 NAND2_1276 (.Y(N5692),.A(N5303),.B(N5304));
NAND2X1 NAND2_1277 (.Y(N5696),.A(N5137),.B(N5305));
NAND2X1 NAND2_1278 (.Y(N5700),.A(N5306),.B(N5140));
NAND2X1 NAND2_1279 (.Y(N5703),.A(N5307),.B(N5308));
NAND2X1 NAND2_1280 (.Y(N5707),.A(N5309),.B(N5310));
NAND2X1 NAND2_1281 (.Y(N5711),.A(N5145),.B(N5311));
AND2X1 AND2_1282 (.Y(N5726),.A(N5166),.B(N4512));
INVX1 NOT1_1283 (.Y(N5727),.A(N5173));
INVX1 NOT1_1284 (.Y(N5728),.A(N5177));
INVX1 NOT1_1285 (.Y(N5730),.A(N5199));
INVX1 NOT1_1286 (.Y(N5731),.A(N5205));
INVX1 NOT1_1287 (.Y(N5732),.A(N5208));
INVX1 NOT1_1288 (.Y(N5733),.A(N5214));
INVX1 NOT1_1289 (.Y(N5734),.A(N5217));
INVX1 NOT1_1290 (.Y(N5735),.A(N5220));
NAND2X1 NAND2_1291 (.Y(N5736),.A(N5365),.B(N5366));
NAND2X1 NAND2_1292 (.Y(N5739),.A(N5363),.B(N5364));
NAND2X1 NAND2_1293 (.Y(N5742),.A(N5369),.B(N5370));
NAND2X1 NAND2_1294 (.Y(N5745),.A(N5367),.B(N5368));
INVX1 NOT1_1295 (.Y(N5755),.A(N5236));
NAND2X1 NAND2_1296 (.Y(N5756),.A(N5332),.B(N5331));
AND2X1 AND2_1297 (.Y(N5954),.A(N5264),.B(N4396));
NAND2X1 NAND2_1298 (.Y(N5955),.A(N1899),.B(N5617));
INVX1 NOT1_1299 (.Y(N5956),.A(N5346));
AND2X1 AND2_1300 (.Y(N6005),.A(N5284),.B(N4456));
AND2X1 AND2_1301 (.Y(N6006),.A(N5284),.B(N4456));
INVX1 NOT1_1302 (.Y(N6023),.A(N5371));
NAND2X1 NAND2_1303 (.Y(N6024),.A(N5371),.B(N5312));
INVX1 NOT1_1304 (.Y(N6025),.A(N5315));
INVX1 NOT1_1305 (.Y(N6028),.A(N5324));
BUFX1 BUFF1_1306 (.Y(N6031),.A(N5319));
BUFX1 BUFF1_1307 (.Y(N6034),.A(N5319));
BUFX1 BUFF1_1308 (.Y(N6037),.A(N5328));
BUFX1 BUFF1_1309 (.Y(N6040),.A(N5328));
INVX1 NOT1_1310 (.Y(N6044),.A(N5385));
OR2X1 OR2_1311 (.Y(N6045),.A(N5166),.B(N5726));
BUFX1 BUFF1_1312 (.Y(N6048),.A(N5264));
BUFX1 BUFF1_1313 (.Y(N6051),.A(N5284));
BUFX1 BUFF1_1314 (.Y(N6054),.A(N5284));
INVX1 NOT1_1315 (.Y(N6065),.A(N5374));
NAND2X1 NAND2_1316 (.Y(N6066),.A(N5374),.B(N5054));
INVX1 NOT1_1317 (.Y(N6067),.A(N5377));
INVX1 NOT1_1318 (.Y(N6068),.A(N5382));
NAND2X1 NAND2_1319 (.Y(N6069),.A(N5382),.B(N5755));
AND2X1 AND2_1320 (.Y(N6071),.A(N5470),.B(N4316));
AND2X1 AND_tmp476 (.Y(ttmp476),.A(N5470),.B(N4320));
AND2X1 AND_tmp477 (.Y(N6072),.A(N5477),.B(ttmp476));
AND2X1 AND_tmp478 (.Y(ttmp478),.A(N4325),.B(N5477));
AND2X1 AND_tmp479 (.Y(ttmp479),.A(N5488),.B(ttmp478));
AND2X1 AND_tmp480 (.Y(N6073),.A(N5470),.B(ttmp479));
AND2X1 AND_tmp481 (.Y(ttmp481),.A(N4385),.B(N4364));
AND2X1 AND_tmp482 (.Y(ttmp482),.A(N5562),.B(ttmp481));
AND2X1 AND_tmp483 (.Y(N6074),.A(N4357),.B(ttmp482));
AND2X1 AND2_1324 (.Y(N6075),.A(N5389),.B(N4280));
AND2X1 AND_tmp484 (.Y(ttmp484),.A(N5389),.B(N4284));
AND2X1 AND_tmp485 (.Y(N6076),.A(N5396),.B(ttmp484));
AND2X1 AND_tmp486 (.Y(ttmp486),.A(N4290),.B(N5396));
AND2X1 AND_tmp487 (.Y(ttmp487),.A(N5407),.B(ttmp486));
AND2X1 AND_tmp488 (.Y(N6077),.A(N5389),.B(ttmp487));
AND2X1 AND_tmp489 (.Y(ttmp489),.A(N4445),.B(N4425));
AND2X1 AND_tmp490 (.Y(ttmp490),.A(N5624),.B(ttmp489));
AND2X1 AND_tmp491 (.Y(N6078),.A(N4418),.B(ttmp490));
INVX1 NOT1_1328 (.Y(N6079),.A(N5418));
AND2X1 AND_tmp492 (.Y(ttmp492),.A(N5407),.B(N5389));
AND2X1 AND_tmp493 (.Y(ttmp493),.A(N5396),.B(ttmp492));
AND2X1 AND_tmp494 (.Y(N6080),.A(N5418),.B(ttmp493));
AND2X1 AND2_1330 (.Y(N6083),.A(N5396),.B(N4284));
AND2X1 AND_tmp495 (.Y(ttmp495),.A(N4290),.B(N5396));
AND2X1 AND_tmp496 (.Y(N6084),.A(N5407),.B(ttmp495));
AND2X1 AND_tmp497 (.Y(ttmp497),.A(N5407),.B(N5396));
AND2X1 AND_tmp498 (.Y(N6085),.A(N5418),.B(ttmp497));
AND2X1 AND2_1333 (.Y(N6086),.A(N5396),.B(N4284));
AND2X1 AND_tmp499 (.Y(ttmp499),.A(N5407),.B(N5396));
AND2X1 AND_tmp500 (.Y(N6087),.A(N4290),.B(ttmp499));
AND2X1 AND2_1335 (.Y(N6088),.A(N5407),.B(N4290));
AND2X1 AND2_1336 (.Y(N6089),.A(N5418),.B(N5407));
AND2X1 AND2_1337 (.Y(N6090),.A(N5407),.B(N4290));
AND2X1 AND_tmp501 (.Y(ttmp501),.A(N5424),.B(N5452));
AND2X1 AND_tmp502 (.Y(ttmp502),.A(N5431),.B(ttmp501));
AND2X1 AND_tmp503 (.Y(ttmp503),.A(N5462),.B(ttmp502));
AND2X1 AND_tmp504 (.Y(N6091),.A(N5441),.B(ttmp503));
AND2X1 AND2_1339 (.Y(N6094),.A(N5424),.B(N4298));
AND2X1 AND_tmp505 (.Y(ttmp505),.A(N5424),.B(N4301));
AND2X1 AND_tmp506 (.Y(N6095),.A(N5431),.B(ttmp505));
AND2X1 AND_tmp507 (.Y(ttmp507),.A(N4305),.B(N5431));
AND2X1 AND_tmp508 (.Y(ttmp508),.A(N5441),.B(ttmp507));
AND2X1 AND_tmp509 (.Y(N6096),.A(N5424),.B(ttmp508));
AND2X1 AND_tmp510 (.Y(ttmp510),.A(N4310),.B(N5431));
AND2X1 AND_tmp511 (.Y(ttmp511),.A(N5452),.B(ttmp510));
AND2X1 AND_tmp512 (.Y(ttmp512),.A(N5441),.B(ttmp511));
AND2X1 AND_tmp513 (.Y(N6097),.A(N5424),.B(ttmp512));
AND2X1 AND2_1343 (.Y(N6098),.A(N5431),.B(N4301));
AND2X1 AND_tmp514 (.Y(ttmp514),.A(N4305),.B(N5431));
AND2X1 AND_tmp515 (.Y(N6099),.A(N5441),.B(ttmp514));
AND2X1 AND_tmp516 (.Y(ttmp516),.A(N4310),.B(N5431));
AND2X1 AND_tmp517 (.Y(ttmp517),.A(N5452),.B(ttmp516));
AND2X1 AND_tmp518 (.Y(N6100),.A(N5441),.B(ttmp517));
AND2X1 AND_tmp519 (.Y(ttmp519),.A(N5452),.B(N5431));
AND2X1 AND_tmp520 (.Y(ttmp520),.A(N4),.B(ttmp519));
AND2X1 AND_tmp521 (.Y(ttmp521),.A(N5462),.B(ttmp520));
AND2X1 AND_tmp522 (.Y(N6101),.A(N5441),.B(ttmp521));
AND2X1 AND2_1347 (.Y(N6102),.A(N4305),.B(N5441));
AND2X1 AND_tmp523 (.Y(ttmp523),.A(N5441),.B(N4310));
AND2X1 AND_tmp524 (.Y(N6103),.A(N5452),.B(ttmp523));
AND2X1 AND_tmp525 (.Y(ttmp525),.A(N5441),.B(N5452));
AND2X1 AND_tmp526 (.Y(ttmp526),.A(N4),.B(ttmp525));
AND2X1 AND_tmp527 (.Y(N6104),.A(N5462),.B(ttmp526));
AND2X1 AND2_1350 (.Y(N6105),.A(N5452),.B(N4310));
AND2X1 AND_tmp528 (.Y(ttmp528),.A(N5462),.B(N5452));
AND2X1 AND_tmp529 (.Y(N6106),.A(N4),.B(ttmp528));
AND2X1 AND2_1352 (.Y(N6107),.A(N4),.B(N5462));
AND2X1 AND_tmp530 (.Y(ttmp530),.A(N5477),.B(N5470));
AND2X1 AND_tmp531 (.Y(ttmp531),.A(N5549),.B(ttmp530));
AND2X1 AND_tmp532 (.Y(N6108),.A(N5488),.B(ttmp531));
AND2X1 AND2_1354 (.Y(N6111),.A(N5477),.B(N4320));
AND2X1 AND_tmp533 (.Y(ttmp533),.A(N4325),.B(N5477));
AND2X1 AND_tmp534 (.Y(N6112),.A(N5488),.B(ttmp533));
AND2X1 AND_tmp535 (.Y(ttmp535),.A(N5488),.B(N5477));
AND2X1 AND_tmp536 (.Y(N6113),.A(N5549),.B(ttmp535));
AND2X1 AND2_1357 (.Y(N6114),.A(N5477),.B(N4320));
AND2X1 AND_tmp537 (.Y(ttmp537),.A(N4325),.B(N5477));
AND2X1 AND_tmp538 (.Y(N6115),.A(N5488),.B(ttmp537));
AND2X1 AND2_1359 (.Y(N6116),.A(N5488),.B(N4325));
AND2X1 AND_tmp539 (.Y(ttmp539),.A(N5506),.B(N5498));
AND2X1 AND_tmp540 (.Y(ttmp540),.A(N5555),.B(ttmp539));
AND2X1 AND_tmp541 (.Y(ttmp541),.A(N5536),.B(ttmp540));
AND2X1 AND_tmp542 (.Y(N6117),.A(N5520),.B(ttmp541));
AND2X1 AND2_1361 (.Y(N6120),.A(N5498),.B(N4332));
AND2X1 AND_tmp543 (.Y(ttmp543),.A(N5498),.B(N4336));
AND2X1 AND_tmp544 (.Y(N6121),.A(N5506),.B(ttmp543));
AND2X1 AND_tmp545 (.Y(ttmp545),.A(N4342),.B(N5506));
AND2X1 AND_tmp546 (.Y(ttmp546),.A(N5520),.B(ttmp545));
AND2X1 AND_tmp547 (.Y(N6122),.A(N5498),.B(ttmp546));
AND2X1 AND_tmp548 (.Y(ttmp548),.A(N4349),.B(N5506));
AND2X1 AND_tmp549 (.Y(ttmp549),.A(N5536),.B(ttmp548));
AND2X1 AND_tmp550 (.Y(ttmp550),.A(N5520),.B(ttmp549));
AND2X1 AND_tmp551 (.Y(N6123),.A(N5498),.B(ttmp550));
AND2X1 AND2_1365 (.Y(N6124),.A(N5506),.B(N4336));
AND2X1 AND_tmp552 (.Y(ttmp552),.A(N4342),.B(N5506));
AND2X1 AND_tmp553 (.Y(N6125),.A(N5520),.B(ttmp552));
AND2X1 AND_tmp554 (.Y(ttmp554),.A(N4349),.B(N5506));
AND2X1 AND_tmp555 (.Y(ttmp555),.A(N5536),.B(ttmp554));
AND2X1 AND_tmp556 (.Y(N6126),.A(N5520),.B(ttmp555));
AND2X1 AND_tmp557 (.Y(ttmp557),.A(N5506),.B(N5536));
AND2X1 AND_tmp558 (.Y(ttmp558),.A(N5555),.B(ttmp557));
AND2X1 AND_tmp559 (.Y(N6127),.A(N5520),.B(ttmp558));
AND2X1 AND2_1369 (.Y(N6128),.A(N5506),.B(N4336));
AND2X1 AND_tmp560 (.Y(ttmp560),.A(N4342),.B(N5506));
AND2X1 AND_tmp561 (.Y(N6129),.A(N5520),.B(ttmp560));
AND2X1 AND_tmp562 (.Y(ttmp562),.A(N4349),.B(N5506));
AND2X1 AND_tmp563 (.Y(ttmp563),.A(N5536),.B(ttmp562));
AND2X1 AND_tmp564 (.Y(N6130),.A(N5520),.B(ttmp563));
AND2X1 AND2_1372 (.Y(N6131),.A(N5520),.B(N4342));
AND2X1 AND_tmp565 (.Y(ttmp565),.A(N5520),.B(N4349));
AND2X1 AND_tmp566 (.Y(N6132),.A(N5536),.B(ttmp565));
AND2X1 AND_tmp567 (.Y(ttmp567),.A(N5520),.B(N5536));
AND2X1 AND_tmp568 (.Y(N6133),.A(N5555),.B(ttmp567));
AND2X1 AND2_1375 (.Y(N6134),.A(N5520),.B(N4342));
AND2X1 AND_tmp569 (.Y(ttmp569),.A(N5520),.B(N4349));
AND2X1 AND_tmp570 (.Y(N6135),.A(N5536),.B(ttmp569));
AND2X1 AND2_1377 (.Y(N6136),.A(N5536),.B(N4349));
AND2X1 AND2_1378 (.Y(N6137),.A(N5549),.B(N5488));
AND2X1 AND2_1379 (.Y(N6138),.A(N5555),.B(N5536));
INVX1 NOT1_1380 (.Y(N6139),.A(N5573));
AND2X1 AND_tmp571 (.Y(ttmp571),.A(N5562),.B(N4357));
AND2X1 AND_tmp572 (.Y(ttmp572),.A(N4364),.B(ttmp571));
AND2X1 AND_tmp573 (.Y(N6140),.A(N5573),.B(ttmp572));
AND2X1 AND_tmp574 (.Y(ttmp574),.A(N4385),.B(N4364));
AND2X1 AND_tmp575 (.Y(N6143),.A(N5562),.B(ttmp574));
AND2X1 AND_tmp576 (.Y(ttmp576),.A(N5562),.B(N4364));
AND2X1 AND_tmp577 (.Y(N6144),.A(N5573),.B(ttmp576));
AND2X1 AND_tmp578 (.Y(ttmp578),.A(N5562),.B(N4364));
AND2X1 AND_tmp579 (.Y(N6145),.A(N4385),.B(ttmp578));
AND2X1 AND2_1385 (.Y(N6146),.A(N5562),.B(N4385));
AND2X1 AND2_1386 (.Y(N6147),.A(N5573),.B(N5562));
AND2X1 AND2_1387 (.Y(N6148),.A(N5562),.B(N4385));
AND2X1 AND_tmp580 (.Y(ttmp580),.A(N5579),.B(N5606));
AND2X1 AND_tmp581 (.Y(ttmp581),.A(N5264),.B(ttmp580));
AND2X1 AND_tmp582 (.Y(ttmp582),.A(N4405),.B(ttmp581));
AND2X1 AND_tmp583 (.Y(N6149),.A(N5595),.B(ttmp582));
AND2X1 AND2_1389 (.Y(N6152),.A(N5579),.B(N4067));
AND2X1 AND_tmp584 (.Y(ttmp584),.A(N5579),.B(N4396));
AND2X1 AND_tmp585 (.Y(N6153),.A(N5264),.B(ttmp584));
AND2X1 AND_tmp586 (.Y(ttmp586),.A(N4400),.B(N5264));
AND2X1 AND_tmp587 (.Y(ttmp587),.A(N5595),.B(ttmp586));
AND2X1 AND_tmp588 (.Y(N6154),.A(N5579),.B(ttmp587));
AND2X1 AND_tmp589 (.Y(ttmp589),.A(N4412),.B(N5264));
AND2X1 AND_tmp590 (.Y(ttmp590),.A(N5606),.B(ttmp589));
AND2X1 AND_tmp591 (.Y(ttmp591),.A(N5595),.B(ttmp590));
AND2X1 AND_tmp592 (.Y(N6155),.A(N5579),.B(ttmp591));
AND2X1 AND_tmp593 (.Y(ttmp593),.A(N4400),.B(N5264));
AND2X1 AND_tmp594 (.Y(N6156),.A(N5595),.B(ttmp593));
AND2X1 AND_tmp595 (.Y(ttmp595),.A(N4412),.B(N5264));
AND2X1 AND_tmp596 (.Y(ttmp596),.A(N5606),.B(ttmp595));
AND2X1 AND_tmp597 (.Y(N6157),.A(N5595),.B(ttmp596));
AND2X1 AND_tmp598 (.Y(ttmp598),.A(N5606),.B(N5264));
AND2X1 AND_tmp599 (.Y(ttmp599),.A(N54),.B(ttmp598));
AND2X1 AND_tmp600 (.Y(ttmp600),.A(N4405),.B(ttmp599));
AND2X1 AND_tmp601 (.Y(N6158),.A(N5595),.B(ttmp600));
AND2X1 AND2_1396 (.Y(N6159),.A(N4400),.B(N5595));
AND2X1 AND_tmp602 (.Y(ttmp602),.A(N5595),.B(N4412));
AND2X1 AND_tmp603 (.Y(N6160),.A(N5606),.B(ttmp602));
AND2X1 AND_tmp604 (.Y(ttmp604),.A(N5595),.B(N5606));
AND2X1 AND_tmp605 (.Y(ttmp605),.A(N54),.B(ttmp604));
AND2X1 AND_tmp606 (.Y(N6161),.A(N4405),.B(ttmp605));
AND2X1 AND2_1399 (.Y(N6162),.A(N5606),.B(N4412));
AND2X1 AND_tmp607 (.Y(ttmp607),.A(N4405),.B(N5606));
AND2X1 AND_tmp608 (.Y(N6163),.A(N54),.B(ttmp607));
NAND2X1 NAND2_1401 (.Y(N6164),.A(N5616),.B(N5955));
AND2X1 AND_tmp609 (.Y(ttmp609),.A(N4425),.B(N4418));
AND2X1 AND_tmp610 (.Y(ttmp610),.A(N5684),.B(ttmp609));
AND2X1 AND_tmp611 (.Y(N6168),.A(N5624),.B(ttmp610));
AND2X1 AND_tmp612 (.Y(ttmp612),.A(N4445),.B(N4425));
AND2X1 AND_tmp613 (.Y(N6171),.A(N5624),.B(ttmp612));
AND2X1 AND_tmp614 (.Y(ttmp614),.A(N5624),.B(N4425));
AND2X1 AND_tmp615 (.Y(N6172),.A(N5684),.B(ttmp614));
AND2X1 AND_tmp616 (.Y(ttmp616),.A(N4445),.B(N4425));
AND2X1 AND_tmp617 (.Y(N6173),.A(N5624),.B(ttmp616));
AND2X1 AND2_1406 (.Y(N6174),.A(N5624),.B(N4445));
AND2X1 AND_tmp618 (.Y(ttmp618),.A(N5284),.B(N5634));
AND2X1 AND_tmp619 (.Y(ttmp619),.A(N4477),.B(ttmp618));
AND2X1 AND_tmp620 (.Y(ttmp620),.A(N5671),.B(ttmp619));
AND2X1 AND_tmp621 (.Y(N6175),.A(N5655),.B(ttmp620));
AND2X1 AND2_1408 (.Y(N6178),.A(N5634),.B(N4080));
AND2X1 AND_tmp622 (.Y(ttmp622),.A(N5634),.B(N4456));
AND2X1 AND_tmp623 (.Y(N6179),.A(N5284),.B(ttmp622));
AND2X1 AND_tmp624 (.Y(ttmp624),.A(N4462),.B(N5284));
AND2X1 AND_tmp625 (.Y(ttmp625),.A(N5655),.B(ttmp624));
AND2X1 AND_tmp626 (.Y(N6180),.A(N5634),.B(ttmp625));
AND2X1 AND_tmp627 (.Y(ttmp627),.A(N4469),.B(N5284));
AND2X1 AND_tmp628 (.Y(ttmp628),.A(N5671),.B(ttmp627));
AND2X1 AND_tmp629 (.Y(ttmp629),.A(N5655),.B(ttmp628));
AND2X1 AND_tmp630 (.Y(N6181),.A(N5634),.B(ttmp629));
AND2X1 AND_tmp631 (.Y(ttmp631),.A(N4462),.B(N5284));
AND2X1 AND_tmp632 (.Y(N6182),.A(N5655),.B(ttmp631));
AND2X1 AND_tmp633 (.Y(ttmp633),.A(N4469),.B(N5284));
AND2X1 AND_tmp634 (.Y(ttmp634),.A(N5671),.B(ttmp633));
AND2X1 AND_tmp635 (.Y(N6183),.A(N5655),.B(ttmp634));
AND2X1 AND_tmp636 (.Y(ttmp636),.A(N5284),.B(N5671));
AND2X1 AND_tmp637 (.Y(ttmp637),.A(N4477),.B(ttmp636));
AND2X1 AND_tmp638 (.Y(N6184),.A(N5655),.B(ttmp637));
AND2X1 AND_tmp639 (.Y(ttmp639),.A(N4462),.B(N5284));
AND2X1 AND_tmp640 (.Y(N6185),.A(N5655),.B(ttmp639));
AND2X1 AND_tmp641 (.Y(ttmp641),.A(N4469),.B(N5284));
AND2X1 AND_tmp642 (.Y(ttmp642),.A(N5671),.B(ttmp641));
AND2X1 AND_tmp643 (.Y(N6186),.A(N5655),.B(ttmp642));
AND2X1 AND2_1417 (.Y(N6187),.A(N5655),.B(N4462));
AND2X1 AND_tmp644 (.Y(ttmp644),.A(N5655),.B(N4469));
AND2X1 AND_tmp645 (.Y(N6188),.A(N5671),.B(ttmp644));
AND2X1 AND_tmp646 (.Y(ttmp646),.A(N5655),.B(N5671));
AND2X1 AND_tmp647 (.Y(N6189),.A(N4477),.B(ttmp646));
AND2X1 AND2_1420 (.Y(N6190),.A(N5655),.B(N4462));
AND2X1 AND_tmp648 (.Y(ttmp648),.A(N5655),.B(N4469));
AND2X1 AND_tmp649 (.Y(N6191),.A(N5671),.B(ttmp648));
AND2X1 AND2_1422 (.Y(N6192),.A(N5671),.B(N4469));
AND2X1 AND2_1423 (.Y(N6193),.A(N5684),.B(N5624));
AND2X1 AND2_1424 (.Y(N6194),.A(N4477),.B(N5671));
INVX1 NOT1_1425 (.Y(N6197),.A(N5692));
INVX1 NOT1_1426 (.Y(N6200),.A(N5696));
INVX1 NOT1_1427 (.Y(N6203),.A(N5703));
INVX1 NOT1_1428 (.Y(N6206),.A(N5707));
BUFX1 BUFF1_1429 (.Y(N6209),.A(N5700));
BUFX1 BUFF1_1430 (.Y(N6212),.A(N5700));
BUFX1 BUFF1_1431 (.Y(N6215),.A(N5711));
BUFX1 BUFF1_1432 (.Y(N6218),.A(N5711));
NAND2X1 NAND2_1433 (.Y(N6221),.A(N5049),.B(N6023));
INVX1 NOT1_1434 (.Y(N6234),.A(N5756));
NAND2X1 NAND2_1435 (.Y(N6235),.A(N5756),.B(N6044));
BUFX1 BUFF1_1436 (.Y(N6238),.A(N5462));
BUFX1 BUFF1_1437 (.Y(N6241),.A(N5389));
BUFX1 BUFF1_1438 (.Y(N6244),.A(N5389));
BUFX1 BUFF1_1439 (.Y(N6247),.A(N5396));
BUFX1 BUFF1_1440 (.Y(N6250),.A(N5396));
BUFX1 BUFF1_1441 (.Y(N6253),.A(N5407));
BUFX1 BUFF1_1442 (.Y(N6256),.A(N5407));
BUFX1 BUFF1_1443 (.Y(N6259),.A(N5424));
BUFX1 BUFF1_1444 (.Y(N6262),.A(N5431));
BUFX1 BUFF1_1445 (.Y(N6265),.A(N5441));
BUFX1 BUFF1_1446 (.Y(N6268),.A(N5452));
BUFX1 BUFF1_1447 (.Y(N6271),.A(N5549));
BUFX1 BUFF1_1448 (.Y(N6274),.A(N5488));
BUFX1 BUFF1_1449 (.Y(N6277),.A(N5470));
BUFX1 BUFF1_1450 (.Y(N6280),.A(N5477));
BUFX1 BUFF1_1451 (.Y(N6283),.A(N5549));
BUFX1 BUFF1_1452 (.Y(N6286),.A(N5488));
BUFX1 BUFF1_1453 (.Y(N6289),.A(N5470));
BUFX1 BUFF1_1454 (.Y(N6292),.A(N5477));
BUFX1 BUFF1_1455 (.Y(N6295),.A(N5555));
BUFX1 BUFF1_1456 (.Y(N6298),.A(N5536));
BUFX1 BUFF1_1457 (.Y(N6301),.A(N5498));
BUFX1 BUFF1_1458 (.Y(N6304),.A(N5520));
BUFX1 BUFF1_1459 (.Y(N6307),.A(N5506));
BUFX1 BUFF1_1460 (.Y(N6310),.A(N5506));
BUFX1 BUFF1_1461 (.Y(N6313),.A(N5555));
BUFX1 BUFF1_1462 (.Y(N6316),.A(N5536));
BUFX1 BUFF1_1463 (.Y(N6319),.A(N5498));
BUFX1 BUFF1_1464 (.Y(N6322),.A(N5520));
BUFX1 BUFF1_1465 (.Y(N6325),.A(N5562));
BUFX1 BUFF1_1466 (.Y(N6328),.A(N5562));
BUFX1 BUFF1_1467 (.Y(N6331),.A(N5579));
BUFX1 BUFF1_1468 (.Y(N6335),.A(N5595));
BUFX1 BUFF1_1469 (.Y(N6338),.A(N5606));
BUFX1 BUFF1_1470 (.Y(N6341),.A(N5684));
BUFX1 BUFF1_1471 (.Y(N6344),.A(N5624));
BUFX1 BUFF1_1472 (.Y(N6347),.A(N5684));
BUFX1 BUFF1_1473 (.Y(N6350),.A(N5624));
BUFX1 BUFF1_1474 (.Y(N6353),.A(N5671));
BUFX1 BUFF1_1475 (.Y(N6356),.A(N5634));
BUFX1 BUFF1_1476 (.Y(N6359),.A(N5655));
BUFX1 BUFF1_1477 (.Y(N6364),.A(N5671));
BUFX1 BUFF1_1478 (.Y(N6367),.A(N5634));
BUFX1 BUFF1_1479 (.Y(N6370),.A(N5655));
INVX1 NOT1_1480 (.Y(N6373),.A(N5736));
INVX1 NOT1_1481 (.Y(N6374),.A(N5739));
INVX1 NOT1_1482 (.Y(N6375),.A(N5742));
INVX1 NOT1_1483 (.Y(N6376),.A(N5745));
NAND2X1 NAND2_1484 (.Y(N6377),.A(N4243),.B(N6065));
NAND2X1 NAND2_1485 (.Y(N6378),.A(N5236),.B(N6068));
OR2X1 OR_tmp650 (.Y(ttmp650),.A(N6072),.B(N6073));
OR2X1 OR_tmp651 (.Y(ttmp651),.A(N4268),.B(ttmp650));
OR2X1 OR_tmp652 (.Y(N6382),.A(N6071),.B(ttmp651));
OR2X1 OR_tmp653 (.Y(ttmp653),.A(N5066),.B(N6074));
OR2X1 OR_tmp654 (.Y(ttmp654),.A(N3968),.B(ttmp653));
OR2X1 OR_tmp655 (.Y(N6386),.A(N5065),.B(ttmp654));
OR2X1 OR_tmp656 (.Y(ttmp656),.A(N6076),.B(N6077));
OR2X1 OR_tmp657 (.Y(ttmp657),.A(N4271),.B(ttmp656));
OR2X1 OR_tmp658 (.Y(N6388),.A(N6075),.B(ttmp657));
OR2X1 OR_tmp659 (.Y(ttmp659),.A(N5068),.B(N6078));
OR2X1 OR_tmp660 (.Y(ttmp660),.A(N3968),.B(ttmp659));
OR2X1 OR_tmp661 (.Y(N6392),.A(N5067),.B(ttmp660));
OR2X1 OR_tmp662 (.Y(ttmp662),.A(N6096),.B(N6097));
OR2X1 OR_tmp663 (.Y(ttmp663),.A(N4297),.B(ttmp662));
OR2X1 OR_tmp664 (.Y(ttmp664),.A(N6094),.B(ttmp663));
OR2X1 OR_tmp665 (.Y(N6397),.A(N6095),.B(ttmp664));
OR2X1 OR2_1491 (.Y(N6411),.A(N4320),.B(N6116));
OR2X1 OR_tmp666 (.Y(ttmp666),.A(N6122),.B(N6123));
OR2X1 OR_tmp667 (.Y(ttmp667),.A(N4331),.B(ttmp666));
OR2X1 OR_tmp668 (.Y(ttmp668),.A(N6120),.B(ttmp667));
OR2X1 OR_tmp669 (.Y(N6415),.A(N6121),.B(ttmp668));
OR2X1 OR2_1493 (.Y(N6419),.A(N4342),.B(N6136));
OR2X1 OR_tmp670 (.Y(ttmp670),.A(N6154),.B(N6155));
OR2X1 OR_tmp671 (.Y(ttmp671),.A(N4392),.B(ttmp670));
OR2X1 OR_tmp672 (.Y(ttmp672),.A(N6152),.B(ttmp671));
OR2X1 OR_tmp673 (.Y(N6427),.A(N6153),.B(ttmp672));
INVX1 NOT1_1495 (.Y(N6434),.A(N6048));
OR2X1 OR2_1496 (.Y(N6437),.A(N4440),.B(N6174));
OR2X1 OR_tmp674 (.Y(ttmp674),.A(N6180),.B(N6181));
OR2X1 OR_tmp675 (.Y(ttmp675),.A(N4451),.B(ttmp674));
OR2X1 OR_tmp676 (.Y(ttmp676),.A(N6178),.B(ttmp675));
OR2X1 OR_tmp677 (.Y(N6441),.A(N6179),.B(ttmp676));
OR2X1 OR2_1498 (.Y(N6445),.A(N4462),.B(N6192));
INVX1 NOT1_1499 (.Y(N6448),.A(N6051));
INVX1 NOT1_1500 (.Y(N6449),.A(N6054));
NAND2X1 NAND2_1501 (.Y(N6466),.A(N6221),.B(N6024));
INVX1 NOT1_1502 (.Y(N6469),.A(N6031));
INVX1 NOT1_1503 (.Y(N6470),.A(N6034));
INVX1 NOT1_1504 (.Y(N6471),.A(N6037));
INVX1 NOT1_1505 (.Y(N6472),.A(N6040));
AND2X1 AND_tmp678 (.Y(ttmp678),.A(N4524),.B(N6031));
AND2X1 AND_tmp679 (.Y(N6473),.A(N5315),.B(ttmp678));
AND2X1 AND_tmp680 (.Y(ttmp680),.A(N5150),.B(N6034));
AND2X1 AND_tmp681 (.Y(N6474),.A(N6025),.B(ttmp680));
AND2X1 AND_tmp682 (.Y(ttmp682),.A(N4532),.B(N6037));
AND2X1 AND_tmp683 (.Y(N6475),.A(N5324),.B(ttmp682));
AND2X1 AND_tmp684 (.Y(ttmp684),.A(N5157),.B(N6040));
AND2X1 AND_tmp685 (.Y(N6476),.A(N6028),.B(ttmp684));
NAND2X1 NAND2_1510 (.Y(N6477),.A(N5385),.B(N6234));
NAND2X1 NAND2_1511 (.Y(N6478),.A(N6045),.B(N132));
OR2X1 OR_tmp686 (.Y(ttmp686),.A(N6084),.B(N6085));
OR2X1 OR_tmp687 (.Y(ttmp687),.A(N4280),.B(ttmp686));
OR2X1 OR_tmp688 (.Y(N6482),.A(N6083),.B(ttmp687));
OR2X1 OR_tmp689 (.Y(ttmp689),.A(N6086),.B(N6087));
NOR2X1 NOR_tmp690 (.Y(N6486),.A(N4280),.B(ttmp689));
OR2X1 OR_tmp691 (.Y(ttmp691),.A(N6088),.B(N6089));
OR2X1 OR_tmp692 (.Y(N6490),.A(N4284),.B(ttmp691));
NOR2X1 NOR2_1515 (.Y(N6494),.A(N4284),.B(N6090));
OR2X1 OR_tmp693 (.Y(ttmp693),.A(N6100),.B(N6101));
OR2X1 OR_tmp694 (.Y(ttmp694),.A(N4298),.B(ttmp693));
OR2X1 OR_tmp695 (.Y(ttmp695),.A(N6098),.B(ttmp694));
OR2X1 OR_tmp696 (.Y(N6500),.A(N6099),.B(ttmp695));
OR2X1 OR_tmp697 (.Y(ttmp697),.A(N6103),.B(N6104));
OR2X1 OR_tmp698 (.Y(ttmp698),.A(N4301),.B(ttmp697));
OR2X1 OR_tmp699 (.Y(N6504),.A(N6102),.B(ttmp698));
OR2X1 OR_tmp700 (.Y(ttmp700),.A(N6105),.B(N6106));
OR2X1 OR_tmp701 (.Y(N6508),.A(N4305),.B(ttmp700));
OR2X1 OR2_1519 (.Y(N6512),.A(N4310),.B(N6107));
OR2X1 OR_tmp702 (.Y(ttmp702),.A(N6112),.B(N6113));
OR2X1 OR_tmp703 (.Y(ttmp703),.A(N4316),.B(ttmp702));
OR2X1 OR_tmp704 (.Y(N6516),.A(N6111),.B(ttmp703));
OR2X1 OR_tmp705 (.Y(ttmp705),.A(N6114),.B(N6115));
NOR2X1 NOR_tmp706 (.Y(N6526),.A(N4316),.B(ttmp705));
OR2X1 OR_tmp707 (.Y(ttmp707),.A(N6132),.B(N6133));
OR2X1 OR_tmp708 (.Y(ttmp708),.A(N4336),.B(ttmp707));
OR2X1 OR_tmp709 (.Y(N6536),.A(N6131),.B(ttmp708));
OR2X1 OR_tmp710 (.Y(ttmp710),.A(N6126),.B(N6127));
OR2X1 OR_tmp711 (.Y(ttmp711),.A(N4332),.B(ttmp710));
OR2X1 OR_tmp712 (.Y(ttmp712),.A(N6124),.B(ttmp711));
OR2X1 OR_tmp713 (.Y(N6539),.A(N6125),.B(ttmp712));
OR2X1 OR_tmp714 (.Y(ttmp714),.A(N6134),.B(N6135));
NOR2X1 NOR_tmp715 (.Y(N6553),.A(N4336),.B(ttmp714));
OR2X1 OR_tmp716 (.Y(ttmp716),.A(N6129),.B(N6130));
OR2X1 OR_tmp717 (.Y(ttmp717),.A(N4332),.B(ttmp716));
NOR2X1 NOR_tmp718 (.Y(N6556),.A(N6128),.B(ttmp717));
OR2X1 OR_tmp719 (.Y(ttmp719),.A(N6143),.B(N6144));
OR2X1 OR_tmp720 (.Y(ttmp720),.A(N4375),.B(ttmp719));
OR2X1 OR_tmp721 (.Y(N6566),.A(N5117),.B(ttmp720));
OR2X1 OR_tmp722 (.Y(ttmp722),.A(N5118),.B(N6145));
NOR2X1 NOR_tmp723 (.Y(N6569),.A(N4375),.B(ttmp722));
OR2X1 OR_tmp724 (.Y(ttmp724),.A(N6146),.B(N6147));
OR2X1 OR_tmp725 (.Y(N6572),.A(N4379),.B(ttmp724));
NOR2X1 NOR2_1529 (.Y(N6575),.A(N4379),.B(N6148));
OR2X1 OR_tmp726 (.Y(ttmp726),.A(N6157),.B(N6158));
OR2X1 OR_tmp727 (.Y(ttmp727),.A(N4067),.B(ttmp726));
OR2X1 OR_tmp728 (.Y(ttmp728),.A(N5954),.B(ttmp727));
OR2X1 OR_tmp729 (.Y(N6580),.A(N6156),.B(ttmp728));
OR2X1 OR_tmp730 (.Y(ttmp730),.A(N6160),.B(N6161));
OR2X1 OR_tmp731 (.Y(ttmp731),.A(N4396),.B(ttmp730));
OR2X1 OR_tmp732 (.Y(N6584),.A(N6159),.B(ttmp731));
OR2X1 OR_tmp733 (.Y(ttmp733),.A(N6162),.B(N6163));
OR2X1 OR_tmp734 (.Y(N6587),.A(N4400),.B(ttmp733));
OR2X1 OR_tmp735 (.Y(ttmp735),.A(N6171),.B(N6172));
OR2X1 OR_tmp736 (.Y(ttmp736),.A(N4436),.B(ttmp735));
OR2X1 OR_tmp737 (.Y(N6592),.A(N5132),.B(ttmp736));
OR2X1 OR_tmp738 (.Y(ttmp738),.A(N5133),.B(N6173));
NOR2X1 NOR_tmp739 (.Y(N6599),.A(N4436),.B(ttmp738));
OR2X1 OR_tmp740 (.Y(ttmp740),.A(N6188),.B(N6189));
OR2X1 OR_tmp741 (.Y(ttmp741),.A(N4456),.B(ttmp740));
OR2X1 OR_tmp742 (.Y(N6606),.A(N6187),.B(ttmp741));
OR2X1 OR_tmp743 (.Y(ttmp743),.A(N6183),.B(N6184));
OR2X1 OR_tmp744 (.Y(ttmp744),.A(N4080),.B(ttmp743));
OR2X1 OR_tmp745 (.Y(ttmp745),.A(N6005),.B(ttmp744));
OR2X1 OR_tmp746 (.Y(N6609),.A(N6182),.B(ttmp745));
OR2X1 OR_tmp747 (.Y(ttmp747),.A(N6190),.B(N6191));
NOR2X1 NOR_tmp748 (.Y(N6619),.A(N4456),.B(ttmp747));
OR2X1 OR_tmp749 (.Y(ttmp749),.A(N6185),.B(N6186));
OR2X1 OR_tmp750 (.Y(ttmp750),.A(N4080),.B(ttmp749));
NOR2X1 NOR_tmp751 (.Y(N6622),.A(N6006),.B(ttmp750));
NAND2X1 NAND2_1539 (.Y(N6630),.A(N5739),.B(N6373));
NAND2X1 NAND2_1540 (.Y(N6631),.A(N5736),.B(N6374));
NAND2X1 NAND2_1541 (.Y(N6632),.A(N5745),.B(N6375));
NAND2X1 NAND2_1542 (.Y(N6633),.A(N5742),.B(N6376));
NAND2X1 NAND2_1543 (.Y(N6634),.A(N6377),.B(N6066));
NAND2X1 NAND2_1544 (.Y(N6637),.A(N6069),.B(N6378));
INVX1 NOT1_1545 (.Y(N6640),.A(N6164));
AND2X1 AND2_1546 (.Y(N6641),.A(N6108),.B(N6117));
AND2X1 AND2_1547 (.Y(N6643),.A(N6140),.B(N6149));
AND2X1 AND2_1548 (.Y(N6646),.A(N6168),.B(N6175));
AND2X1 AND2_1549 (.Y(N6648),.A(N6080),.B(N6091));
NAND2X1 NAND2_1550 (.Y(N6650),.A(N6238),.B(N2637));
INVX1 NOT1_1551 (.Y(N6651),.A(N6238));
INVX1 NOT1_1552 (.Y(N6653),.A(N6241));
INVX1 NOT1_1553 (.Y(N6655),.A(N6244));
INVX1 NOT1_1554 (.Y(N6657),.A(N6247));
INVX1 NOT1_1555 (.Y(N6659),.A(N6250));
NAND2X1 NAND2_1556 (.Y(N6660),.A(N6253),.B(N5087));
INVX1 NOT1_1557 (.Y(N6661),.A(N6253));
NAND2X1 NAND2_1558 (.Y(N6662),.A(N6256),.B(N5469));
INVX1 NOT1_1559 (.Y(N6663),.A(N6256));
AND2X1 AND2_1560 (.Y(N6664),.A(N6091),.B(N4));
INVX1 NOT1_1561 (.Y(N6666),.A(N6259));
INVX1 NOT1_1562 (.Y(N6668),.A(N6262));
INVX1 NOT1_1563 (.Y(N6670),.A(N6265));
INVX1 NOT1_1564 (.Y(N6672),.A(N6268));
INVX1 NOT1_1565 (.Y(N6675),.A(N6117));
INVX1 NOT1_1566 (.Y(N6680),.A(N6280));
INVX1 NOT1_1567 (.Y(N6681),.A(N6292));
INVX1 NOT1_1568 (.Y(N6682),.A(N6307));
INVX1 NOT1_1569 (.Y(N6683),.A(N6310));
NAND2X1 NAND2_1570 (.Y(N6689),.A(N6325),.B(N5120));
INVX1 NOT1_1571 (.Y(N6690),.A(N6325));
NAND2X1 NAND2_1572 (.Y(N6691),.A(N6328),.B(N5622));
INVX1 NOT1_1573 (.Y(N6692),.A(N6328));
AND2X1 AND2_1574 (.Y(N6693),.A(N6149),.B(N54));
INVX1 NOT1_1575 (.Y(N6695),.A(N6331));
INVX1 NOT1_1576 (.Y(N6698),.A(N6335));
NAND2X1 NAND2_1577 (.Y(N6699),.A(N6338),.B(N5956));
INVX1 NOT1_1578 (.Y(N6700),.A(N6338));
INVX1 NOT1_1579 (.Y(N6703),.A(N6175));
INVX1 NOT1_1580 (.Y(N6708),.A(N6209));
INVX1 NOT1_1581 (.Y(N6709),.A(N6212));
INVX1 NOT1_1582 (.Y(N6710),.A(N6215));
INVX1 NOT1_1583 (.Y(N6711),.A(N6218));
AND2X1 AND_tmp752 (.Y(ttmp752),.A(N5692),.B(N6209));
AND2X1 AND_tmp753 (.Y(N6712),.A(N5696),.B(ttmp752));
AND2X1 AND_tmp754 (.Y(ttmp754),.A(N6197),.B(N6212));
AND2X1 AND_tmp755 (.Y(N6713),.A(N6200),.B(ttmp754));
AND2X1 AND_tmp756 (.Y(ttmp756),.A(N5703),.B(N6215));
AND2X1 AND_tmp757 (.Y(N6714),.A(N5707),.B(ttmp756));
AND2X1 AND_tmp758 (.Y(ttmp758),.A(N6203),.B(N6218));
AND2X1 AND_tmp759 (.Y(N6715),.A(N6206),.B(ttmp758));
BUFX1 BUFF1_1588 (.Y(N6716),.A(N6466));
AND2X1 AND_tmp760 (.Y(ttmp760),.A(N1777),.B(N3130));
AND2X1 AND_tmp761 (.Y(N6718),.A(N6164),.B(ttmp760));
AND2X1 AND_tmp762 (.Y(ttmp762),.A(N5315),.B(N6469));
AND2X1 AND_tmp763 (.Y(N6719),.A(N5150),.B(ttmp762));
AND2X1 AND_tmp764 (.Y(ttmp764),.A(N6025),.B(N6470));
AND2X1 AND_tmp765 (.Y(N6720),.A(N4524),.B(ttmp764));
AND2X1 AND_tmp766 (.Y(ttmp766),.A(N5324),.B(N6471));
AND2X1 AND_tmp767 (.Y(N6721),.A(N5157),.B(ttmp766));
AND2X1 AND_tmp768 (.Y(ttmp768),.A(N6028),.B(N6472));
AND2X1 AND_tmp769 (.Y(N6722),.A(N4532),.B(ttmp768));
NAND2X1 NAND2_1594 (.Y(N6724),.A(N6477),.B(N6235));
INVX1 NOT1_1595 (.Y(N6739),.A(N6271));
INVX1 NOT1_1596 (.Y(N6740),.A(N6274));
INVX1 NOT1_1597 (.Y(N6741),.A(N6277));
INVX1 NOT1_1598 (.Y(N6744),.A(N6283));
INVX1 NOT1_1599 (.Y(N6745),.A(N6286));
INVX1 NOT1_1600 (.Y(N6746),.A(N6289));
INVX1 NOT1_1601 (.Y(N6751),.A(N6295));
INVX1 NOT1_1602 (.Y(N6752),.A(N6298));
INVX1 NOT1_1603 (.Y(N6753),.A(N6301));
INVX1 NOT1_1604 (.Y(N6754),.A(N6304));
INVX1 NOT1_1605 (.Y(N6755),.A(N6322));
INVX1 NOT1_1606 (.Y(N6760),.A(N6313));
INVX1 NOT1_1607 (.Y(N6761),.A(N6316));
INVX1 NOT1_1608 (.Y(N6762),.A(N6319));
INVX1 NOT1_1609 (.Y(N6772),.A(N6341));
INVX1 NOT1_1610 (.Y(N6773),.A(N6344));
INVX1 NOT1_1611 (.Y(N6776),.A(N6347));
INVX1 NOT1_1612 (.Y(N6777),.A(N6350));
INVX1 NOT1_1613 (.Y(N6782),.A(N6353));
INVX1 NOT1_1614 (.Y(N6783),.A(N6356));
INVX1 NOT1_1615 (.Y(N6784),.A(N6359));
INVX1 NOT1_1616 (.Y(N6785),.A(N6370));
INVX1 NOT1_1617 (.Y(N6790),.A(N6364));
INVX1 NOT1_1618 (.Y(N6791),.A(N6367));
NAND2X1 NAND2_1619 (.Y(N6792),.A(N6630),.B(N6631));
NAND2X1 NAND2_1620 (.Y(N6795),.A(N6632),.B(N6633));
AND2X1 AND2_1621 (.Y(N6801),.A(N6108),.B(N6415));
AND2X1 AND2_1622 (.Y(N6802),.A(N6427),.B(N6140));
AND2X1 AND2_1623 (.Y(N6803),.A(N6397),.B(N6080));
AND2X1 AND2_1624 (.Y(N6804),.A(N6168),.B(N6441));
INVX1 NOT1_1625 (.Y(N6805),.A(N6466));
NAND2X1 NAND2_1626 (.Y(N6806),.A(N1851),.B(N6651));
INVX1 NOT1_1627 (.Y(N6807),.A(N6482));
NAND2X1 NAND2_1628 (.Y(N6808),.A(N6482),.B(N6653));
INVX1 NOT1_1629 (.Y(N6809),.A(N6486));
NAND2X1 NAND2_1630 (.Y(N6810),.A(N6486),.B(N6655));
INVX1 NOT1_1631 (.Y(N6811),.A(N6490));
NAND2X1 NAND2_1632 (.Y(N6812),.A(N6490),.B(N6657));
INVX1 NOT1_1633 (.Y(N6813),.A(N6494));
NAND2X1 NAND2_1634 (.Y(N6814),.A(N6494),.B(N6659));
NAND2X1 NAND2_1635 (.Y(N6815),.A(N4575),.B(N6661));
NAND2X1 NAND2_1636 (.Y(N6816),.A(N5169),.B(N6663));
OR2X1 OR2_1637 (.Y(N6817),.A(N6397),.B(N6664));
INVX1 NOT1_1638 (.Y(N6823),.A(N6500));
NAND2X1 NAND2_1639 (.Y(N6824),.A(N6500),.B(N6666));
INVX1 NOT1_1640 (.Y(N6825),.A(N6504));
NAND2X1 NAND2_1641 (.Y(N6826),.A(N6504),.B(N6668));
INVX1 NOT1_1642 (.Y(N6827),.A(N6508));
NAND2X1 NAND2_1643 (.Y(N6828),.A(N6508),.B(N6670));
INVX1 NOT1_1644 (.Y(N6829),.A(N6512));
NAND2X1 NAND2_1645 (.Y(N6830),.A(N6512),.B(N6672));
INVX1 NOT1_1646 (.Y(N6831),.A(N6415));
INVX1 NOT1_1647 (.Y(N6834),.A(N6566));
NAND2X1 NAND2_1648 (.Y(N6835),.A(N6566),.B(N5618));
INVX1 NOT1_1649 (.Y(N6836),.A(N6569));
NAND2X1 NAND2_1650 (.Y(N6837),.A(N6569),.B(N5619));
INVX1 NOT1_1651 (.Y(N6838),.A(N6572));
NAND2X1 NAND2_1652 (.Y(N6839),.A(N6572),.B(N5620));
INVX1 NOT1_1653 (.Y(N6840),.A(N6575));
NAND2X1 NAND2_1654 (.Y(N6841),.A(N6575),.B(N5621));
NAND2X1 NAND2_1655 (.Y(N6842),.A(N4627),.B(N6690));
NAND2X1 NAND2_1656 (.Y(N6843),.A(N5195),.B(N6692));
OR2X1 OR2_1657 (.Y(N6844),.A(N6427),.B(N6693));
INVX1 NOT1_1658 (.Y(N6850),.A(N6580));
NAND2X1 NAND2_1659 (.Y(N6851),.A(N6580),.B(N6695));
INVX1 NOT1_1660 (.Y(N6852),.A(N6584));
NAND2X1 NAND2_1661 (.Y(N6853),.A(N6584),.B(N6434));
INVX1 NOT1_1662 (.Y(N6854),.A(N6587));
NAND2X1 NAND2_1663 (.Y(N6855),.A(N6587),.B(N6698));
NAND2X1 NAND2_1664 (.Y(N6856),.A(N5346),.B(N6700));
INVX1 NOT1_1665 (.Y(N6857),.A(N6441));
AND2X1 AND_tmp770 (.Y(ttmp770),.A(N5696),.B(N6708));
AND2X1 AND_tmp771 (.Y(N6860),.A(N6197),.B(ttmp770));
AND2X1 AND_tmp772 (.Y(ttmp772),.A(N6200),.B(N6709));
AND2X1 AND_tmp773 (.Y(N6861),.A(N5692),.B(ttmp772));
AND2X1 AND_tmp774 (.Y(ttmp774),.A(N5707),.B(N6710));
AND2X1 AND_tmp775 (.Y(N6862),.A(N6203),.B(ttmp774));
AND2X1 AND_tmp776 (.Y(ttmp776),.A(N6206),.B(N6711));
AND2X1 AND_tmp777 (.Y(N6863),.A(N5703),.B(ttmp776));
OR2X1 OR_tmp778 (.Y(ttmp778),.A(N6718),.B(N3785));
OR2X1 OR_tmp779 (.Y(N6866),.A(N4197),.B(ttmp778));
NOR2X1 NOR2_1671 (.Y(N6872),.A(N6719),.B(N6473));
NOR2X1 NOR2_1672 (.Y(N6873),.A(N6720),.B(N6474));
NOR2X1 NOR2_1673 (.Y(N6874),.A(N6721),.B(N6475));
NOR2X1 NOR2_1674 (.Y(N6875),.A(N6722),.B(N6476));
INVX1 NOT1_1675 (.Y(N6876),.A(N6637));
BUFX1 BUFF1_1676 (.Y(N6877),.A(N6724));
AND2X1 AND2_1677 (.Y(N6879),.A(N6045),.B(N6478));
AND2X1 AND2_1678 (.Y(N6880),.A(N6478),.B(N132));
OR2X1 OR2_1679 (.Y(N6881),.A(N6411),.B(N6137));
INVX1 NOT1_1680 (.Y(N6884),.A(N6516));
INVX1 NOT1_1681 (.Y(N6885),.A(N6411));
INVX1 NOT1_1682 (.Y(N6888),.A(N6526));
INVX1 NOT1_1683 (.Y(N6889),.A(N6536));
NAND2X1 NAND2_1684 (.Y(N6890),.A(N6536),.B(N5176));
OR2X1 OR2_1685 (.Y(N6891),.A(N6419),.B(N6138));
INVX1 NOT1_1686 (.Y(N6894),.A(N6539));
INVX1 NOT1_1687 (.Y(N6895),.A(N6553));
NAND2X1 NAND2_1688 (.Y(N6896),.A(N6553),.B(N5728));
INVX1 NOT1_1689 (.Y(N6897),.A(N6419));
INVX1 NOT1_1690 (.Y(N6900),.A(N6556));
OR2X1 OR2_1691 (.Y(N6901),.A(N6437),.B(N6193));
INVX1 NOT1_1692 (.Y(N6904),.A(N6592));
INVX1 NOT1_1693 (.Y(N6905),.A(N6437));
INVX1 NOT1_1694 (.Y(N6908),.A(N6599));
OR2X1 OR2_1695 (.Y(N6909),.A(N6445),.B(N6194));
INVX1 NOT1_1696 (.Y(N6912),.A(N6606));
INVX1 NOT1_1697 (.Y(N6913),.A(N6609));
INVX1 NOT1_1698 (.Y(N6914),.A(N6619));
NAND2X1 NAND2_1699 (.Y(N6915),.A(N6619),.B(N5734));
INVX1 NOT1_1700 (.Y(N6916),.A(N6445));
INVX1 NOT1_1701 (.Y(N6919),.A(N6622));
INVX1 NOT1_1702 (.Y(N6922),.A(N6634));
NAND2X1 NAND2_1703 (.Y(N6923),.A(N6634),.B(N6067));
OR2X1 OR2_1704 (.Y(N6924),.A(N6382),.B(N6801));
OR2X1 OR2_1705 (.Y(N6925),.A(N6386),.B(N6802));
OR2X1 OR2_1706 (.Y(N6926),.A(N6388),.B(N6803));
OR2X1 OR2_1707 (.Y(N6927),.A(N6392),.B(N6804));
INVX1 NOT1_1708 (.Y(N6930),.A(N6724));
NAND2X1 NAND2_1709 (.Y(N6932),.A(N6650),.B(N6806));
NAND2X1 NAND2_1710 (.Y(N6935),.A(N6241),.B(N6807));
NAND2X1 NAND2_1711 (.Y(N6936),.A(N6244),.B(N6809));
NAND2X1 NAND2_1712 (.Y(N6937),.A(N6247),.B(N6811));
NAND2X1 NAND2_1713 (.Y(N6938),.A(N6250),.B(N6813));
NAND2X1 NAND2_1714 (.Y(N6939),.A(N6660),.B(N6815));
NAND2X1 NAND2_1715 (.Y(N6940),.A(N6662),.B(N6816));
NAND2X1 NAND2_1716 (.Y(N6946),.A(N6259),.B(N6823));
NAND2X1 NAND2_1717 (.Y(N6947),.A(N6262),.B(N6825));
NAND2X1 NAND2_1718 (.Y(N6948),.A(N6265),.B(N6827));
NAND2X1 NAND2_1719 (.Y(N6949),.A(N6268),.B(N6829));
NAND2X1 NAND2_1720 (.Y(N6953),.A(N5183),.B(N6834));
NAND2X1 NAND2_1721 (.Y(N6954),.A(N5186),.B(N6836));
NAND2X1 NAND2_1722 (.Y(N6955),.A(N5189),.B(N6838));
NAND2X1 NAND2_1723 (.Y(N6956),.A(N5192),.B(N6840));
NAND2X1 NAND2_1724 (.Y(N6957),.A(N6689),.B(N6842));
NAND2X1 NAND2_1725 (.Y(N6958),.A(N6691),.B(N6843));
NAND2X1 NAND2_1726 (.Y(N6964),.A(N6331),.B(N6850));
NAND2X1 NAND2_1727 (.Y(N6965),.A(N6048),.B(N6852));
NAND2X1 NAND2_1728 (.Y(N6966),.A(N6335),.B(N6854));
NAND2X1 NAND2_1729 (.Y(N6967),.A(N6699),.B(N6856));
NOR2X1 NOR2_1730 (.Y(N6973),.A(N6860),.B(N6712));
NOR2X1 NOR2_1731 (.Y(N6974),.A(N6861),.B(N6713));
NOR2X1 NOR2_1732 (.Y(N6975),.A(N6862),.B(N6714));
NOR2X1 NOR2_1733 (.Y(N6976),.A(N6863),.B(N6715));
INVX1 NOT1_1734 (.Y(N6977),.A(N6792));
INVX1 NOT1_1735 (.Y(N6978),.A(N6795));
OR2X1 OR2_1736 (.Y(N6979),.A(N6879),.B(N6880));
NAND2X1 NAND2_1737 (.Y(N6987),.A(N4608),.B(N6889));
NAND2X1 NAND2_1738 (.Y(N6990),.A(N5177),.B(N6895));
NAND2X1 NAND2_1739 (.Y(N6999),.A(N5217),.B(N6914));
NAND2X1 NAND2_1740 (.Y(N7002),.A(N5377),.B(N6922));
NAND2X1 NAND2_1741 (.Y(N7003),.A(N6873),.B(N6872));
NAND2X1 NAND2_1742 (.Y(N7006),.A(N6875),.B(N6874));
AND2X1 AND_tmp780 (.Y(ttmp780),.A(N2681),.B(N2692));
AND2X1 AND_tmp781 (.Y(N7011),.A(N6866),.B(ttmp780));
AND2X1 AND_tmp782 (.Y(ttmp782),.A(N2756),.B(N2767));
AND2X1 AND_tmp783 (.Y(N7012),.A(N6866),.B(ttmp782));
AND2X1 AND_tmp784 (.Y(ttmp784),.A(N2779),.B(N2790));
AND2X1 AND_tmp785 (.Y(N7013),.A(N6866),.B(ttmp784));
INVX1 NOT1_1746 (.Y(N7015),.A(N6866));
AND2X1 AND_tmp786 (.Y(ttmp786),.A(N2801),.B(N2812));
AND2X1 AND_tmp787 (.Y(N7016),.A(N6866),.B(ttmp786));
NAND2X1 NAND2_1748 (.Y(N7018),.A(N6935),.B(N6808));
NAND2X1 NAND2_1749 (.Y(N7019),.A(N6936),.B(N6810));
NAND2X1 NAND2_1750 (.Y(N7020),.A(N6937),.B(N6812));
NAND2X1 NAND2_1751 (.Y(N7021),.A(N6938),.B(N6814));
INVX1 NOT1_1752 (.Y(N7022),.A(N6939));
INVX1 NOT1_1753 (.Y(N7023),.A(N6817));
NAND2X1 NAND2_1754 (.Y(N7028),.A(N6946),.B(N6824));
NAND2X1 NAND2_1755 (.Y(N7031),.A(N6947),.B(N6826));
NAND2X1 NAND2_1756 (.Y(N7034),.A(N6948),.B(N6828));
NAND2X1 NAND2_1757 (.Y(N7037),.A(N6949),.B(N6830));
AND2X1 AND2_1758 (.Y(N7040),.A(N6817),.B(N6079));
AND2X1 AND2_1759 (.Y(N7041),.A(N6831),.B(N6675));
NAND2X1 NAND2_1760 (.Y(N7044),.A(N6953),.B(N6835));
NAND2X1 NAND2_1761 (.Y(N7045),.A(N6954),.B(N6837));
NAND2X1 NAND2_1762 (.Y(N7046),.A(N6955),.B(N6839));
NAND2X1 NAND2_1763 (.Y(N7047),.A(N6956),.B(N6841));
INVX1 NOT1_1764 (.Y(N7048),.A(N6957));
INVX1 NOT1_1765 (.Y(N7049),.A(N6844));
NAND2X1 NAND2_1766 (.Y(N7054),.A(N6964),.B(N6851));
NAND2X1 NAND2_1767 (.Y(N7057),.A(N6965),.B(N6853));
NAND2X1 NAND2_1768 (.Y(N7060),.A(N6966),.B(N6855));
AND2X1 AND2_1769 (.Y(N7064),.A(N6844),.B(N6139));
AND2X1 AND2_1770 (.Y(N7065),.A(N6857),.B(N6703));
INVX1 NOT1_1771 (.Y(N7072),.A(N6881));
NAND2X1 NAND2_1772 (.Y(N7073),.A(N6881),.B(N5172));
INVX1 NOT1_1773 (.Y(N7074),.A(N6885));
NAND2X1 NAND2_1774 (.Y(N7075),.A(N6885),.B(N5727));
NAND2X1 NAND2_1775 (.Y(N7076),.A(N6890),.B(N6987));
INVX1 NOT1_1776 (.Y(N7079),.A(N6891));
NAND2X1 NAND2_1777 (.Y(N7080),.A(N6896),.B(N6990));
INVX1 NOT1_1778 (.Y(N7083),.A(N6897));
INVX1 NOT1_1779 (.Y(N7084),.A(N6901));
NAND2X1 NAND2_1780 (.Y(N7085),.A(N6901),.B(N5198));
INVX1 NOT1_1781 (.Y(N7086),.A(N6905));
NAND2X1 NAND2_1782 (.Y(N7087),.A(N6905),.B(N5731));
INVX1 NOT1_1783 (.Y(N7088),.A(N6909));
NAND2X1 NAND2_1784 (.Y(N7089),.A(N6909),.B(N6912));
NAND2X1 NAND2_1785 (.Y(N7090),.A(N6915),.B(N6999));
INVX1 NOT1_1786 (.Y(N7093),.A(N6916));
NAND2X1 NAND2_1787 (.Y(N7094),.A(N6974),.B(N6973));
NAND2X1 NAND2_1788 (.Y(N7097),.A(N6976),.B(N6975));
NAND2X1 NAND2_1789 (.Y(N7101),.A(N7002),.B(N6923));
INVX1 NOT1_1790 (.Y(N7105),.A(N6932));
INVX1 NOT1_1791 (.Y(N7110),.A(N6967));
AND2X1 AND_tmp788 (.Y(ttmp788),.A(N603),.B(N1755));
AND2X1 AND_tmp789 (.Y(N7114),.A(N6979),.B(ttmp788));
INVX1 NOT1_1793 (.Y(N7115),.A(N7019));
INVX1 NOT1_1794 (.Y(N7116),.A(N7021));
AND2X1 AND2_1795 (.Y(N7125),.A(N6817),.B(N7018));
AND2X1 AND2_1796 (.Y(N7126),.A(N6817),.B(N7020));
AND2X1 AND2_1797 (.Y(N7127),.A(N6817),.B(N7022));
INVX1 NOT1_1798 (.Y(N7130),.A(N7045));
INVX1 NOT1_1799 (.Y(N7131),.A(N7047));
AND2X1 AND2_1800 (.Y(N7139),.A(N6844),.B(N7044));
AND2X1 AND2_1801 (.Y(N7140),.A(N6844),.B(N7046));
AND2X1 AND2_1802 (.Y(N7141),.A(N6844),.B(N7048));
AND2X1 AND_tmp790 (.Y(ttmp790),.A(N1761),.B(N3108));
AND2X1 AND_tmp791 (.Y(N7146),.A(N6932),.B(ttmp790));
AND2X1 AND_tmp792 (.Y(ttmp792),.A(N1777),.B(N3130));
AND2X1 AND_tmp793 (.Y(N7147),.A(N6967),.B(ttmp792));
INVX1 NOT1_1805 (.Y(N7149),.A(N7003));
INVX1 NOT1_1806 (.Y(N7150),.A(N7006));
NAND2X1 NAND2_1807 (.Y(N7151),.A(N7006),.B(N6876));
NAND2X1 NAND2_1808 (.Y(N7152),.A(N4605),.B(N7072));
NAND2X1 NAND2_1809 (.Y(N7153),.A(N5173),.B(N7074));
NAND2X1 NAND2_1810 (.Y(N7158),.A(N4646),.B(N7084));
NAND2X1 NAND2_1811 (.Y(N7159),.A(N5205),.B(N7086));
NAND2X1 NAND2_1812 (.Y(N7160),.A(N6606),.B(N7088));
INVX1 NOT1_1813 (.Y(N7166),.A(N7037));
INVX1 NOT1_1814 (.Y(N7167),.A(N7034));
INVX1 NOT1_1815 (.Y(N7168),.A(N7031));
INVX1 NOT1_1816 (.Y(N7169),.A(N7028));
INVX1 NOT1_1817 (.Y(N7170),.A(N7060));
INVX1 NOT1_1818 (.Y(N7171),.A(N7057));
INVX1 NOT1_1819 (.Y(N7172),.A(N7054));
AND2X1 AND2_1820 (.Y(N7173),.A(N7115),.B(N7023));
AND2X1 AND2_1821 (.Y(N7174),.A(N7116),.B(N7023));
AND2X1 AND2_1822 (.Y(N7175),.A(N6940),.B(N7023));
AND2X1 AND2_1823 (.Y(N7176),.A(N5418),.B(N7023));
INVX1 NOT1_1824 (.Y(N7177),.A(N7041));
AND2X1 AND2_1825 (.Y(N7178),.A(N7130),.B(N7049));
AND2X1 AND2_1826 (.Y(N7179),.A(N7131),.B(N7049));
AND2X1 AND2_1827 (.Y(N7180),.A(N6958),.B(N7049));
AND2X1 AND2_1828 (.Y(N7181),.A(N5573),.B(N7049));
INVX1 NOT1_1829 (.Y(N7182),.A(N7065));
INVX1 NOT1_1830 (.Y(N7183),.A(N7094));
NAND2X1 NAND2_1831 (.Y(N7184),.A(N7094),.B(N6977));
INVX1 NOT1_1832 (.Y(N7185),.A(N7097));
NAND2X1 NAND2_1833 (.Y(N7186),.A(N7097),.B(N6978));
AND2X1 AND_tmp794 (.Y(ttmp794),.A(N1761),.B(N3108));
AND2X1 AND_tmp795 (.Y(N7187),.A(N7037),.B(ttmp794));
AND2X1 AND_tmp796 (.Y(ttmp796),.A(N1761),.B(N3108));
AND2X1 AND_tmp797 (.Y(N7188),.A(N7034),.B(ttmp796));
AND2X1 AND_tmp798 (.Y(ttmp798),.A(N1761),.B(N3108));
AND2X1 AND_tmp799 (.Y(N7189),.A(N7031),.B(ttmp798));
OR2X1 OR_tmp800 (.Y(ttmp800),.A(N7146),.B(N3781));
OR2X1 OR_tmp801 (.Y(N7190),.A(N4956),.B(ttmp800));
AND2X1 AND_tmp802 (.Y(ttmp802),.A(N1777),.B(N3130));
AND2X1 AND_tmp803 (.Y(N7196),.A(N7060),.B(ttmp802));
AND2X1 AND_tmp804 (.Y(ttmp804),.A(N1777),.B(N3130));
AND2X1 AND_tmp805 (.Y(N7197),.A(N7057),.B(ttmp804));
OR2X1 OR_tmp806 (.Y(ttmp806),.A(N7147),.B(N3786));
OR2X1 OR_tmp807 (.Y(N7198),.A(N4960),.B(ttmp806));
NAND2X1 NAND2_1841 (.Y(N7204),.A(N7101),.B(N7149));
INVX1 NOT1_1842 (.Y(N7205),.A(N7101));
NAND2X1 NAND2_1843 (.Y(N7206),.A(N6637),.B(N7150));
AND2X1 AND_tmp808 (.Y(ttmp808),.A(N1793),.B(N3158));
AND2X1 AND_tmp809 (.Y(N7207),.A(N7028),.B(ttmp808));
AND2X1 AND_tmp810 (.Y(ttmp810),.A(N1807),.B(N3180));
AND2X1 AND_tmp811 (.Y(N7208),.A(N7054),.B(ttmp810));
NAND2X1 NAND2_1846 (.Y(N7209),.A(N7073),.B(N7152));
NAND2X1 NAND2_1847 (.Y(N7212),.A(N7075),.B(N7153));
INVX1 NOT1_1848 (.Y(N7215),.A(N7076));
NAND2X1 NAND2_1849 (.Y(N7216),.A(N7076),.B(N7079));
INVX1 NOT1_1850 (.Y(N7217),.A(N7080));
NAND2X1 NAND2_1851 (.Y(N7218),.A(N7080),.B(N7083));
NAND2X1 NAND2_1852 (.Y(N7219),.A(N7085),.B(N7158));
NAND2X1 NAND2_1853 (.Y(N7222),.A(N7087),.B(N7159));
NAND2X1 NAND2_1854 (.Y(N7225),.A(N7089),.B(N7160));
INVX1 NOT1_1855 (.Y(N7228),.A(N7090));
NAND2X1 NAND2_1856 (.Y(N7229),.A(N7090),.B(N7093));
OR2X1 OR2_1857 (.Y(N7236),.A(N7173),.B(N7125));
OR2X1 OR2_1858 (.Y(N7239),.A(N7174),.B(N7126));
OR2X1 OR2_1859 (.Y(N7242),.A(N7175),.B(N7127));
OR2X1 OR2_1860 (.Y(N7245),.A(N7176),.B(N7040));
OR2X1 OR2_1861 (.Y(N7250),.A(N7178),.B(N7139));
OR2X1 OR2_1862 (.Y(N7257),.A(N7179),.B(N7140));
OR2X1 OR2_1863 (.Y(N7260),.A(N7180),.B(N7141));
OR2X1 OR2_1864 (.Y(N7263),.A(N7181),.B(N7064));
NAND2X1 NAND2_1865 (.Y(N7268),.A(N6792),.B(N7183));
NAND2X1 NAND2_1866 (.Y(N7269),.A(N6795),.B(N7185));
OR2X1 OR_tmp812 (.Y(ttmp812),.A(N7187),.B(N3782));
OR2X1 OR_tmp813 (.Y(N7270),.A(N4957),.B(ttmp812));
OR2X1 OR_tmp814 (.Y(ttmp814),.A(N7188),.B(N3783));
OR2X1 OR_tmp815 (.Y(N7276),.A(N4958),.B(ttmp814));
OR2X1 OR_tmp816 (.Y(ttmp816),.A(N7189),.B(N3784));
OR2X1 OR_tmp817 (.Y(N7282),.A(N4959),.B(ttmp816));
OR2X1 OR_tmp818 (.Y(ttmp818),.A(N7196),.B(N3787));
OR2X1 OR_tmp819 (.Y(N7288),.A(N4961),.B(ttmp818));
OR2X1 OR_tmp820 (.Y(ttmp820),.A(N7197),.B(N3788));
OR2X1 OR_tmp821 (.Y(N7294),.A(N3998),.B(ttmp820));
NAND2X1 NAND2_1872 (.Y(N7300),.A(N7003),.B(N7205));
NAND2X1 NAND2_1873 (.Y(N7301),.A(N7206),.B(N7151));
OR2X1 OR_tmp822 (.Y(ttmp822),.A(N7207),.B(N3800));
OR2X1 OR_tmp823 (.Y(N7304),.A(N4980),.B(ttmp822));
OR2X1 OR_tmp824 (.Y(ttmp824),.A(N7208),.B(N3805));
OR2X1 OR_tmp825 (.Y(N7310),.A(N4984),.B(ttmp824));
NAND2X1 NAND2_1876 (.Y(N7320),.A(N6891),.B(N7215));
NAND2X1 NAND2_1877 (.Y(N7321),.A(N6897),.B(N7217));
NAND2X1 NAND2_1878 (.Y(N7328),.A(N6916),.B(N7228));
AND2X1 AND_tmp826 (.Y(ttmp826),.A(N1185),.B(N2692));
AND2X1 AND_tmp827 (.Y(N7338),.A(N7190),.B(ttmp826));
AND2X1 AND_tmp828 (.Y(ttmp828),.A(N2681),.B(N2692));
AND2X1 AND_tmp829 (.Y(N7339),.A(N7198),.B(ttmp828));
AND2X1 AND_tmp830 (.Y(ttmp830),.A(N1247),.B(N2767));
AND2X1 AND_tmp831 (.Y(N7340),.A(N7190),.B(ttmp830));
AND2X1 AND_tmp832 (.Y(ttmp832),.A(N2756),.B(N2767));
AND2X1 AND_tmp833 (.Y(N7341),.A(N7198),.B(ttmp832));
AND2X1 AND_tmp834 (.Y(ttmp834),.A(N1327),.B(N2790));
AND2X1 AND_tmp835 (.Y(N7342),.A(N7190),.B(ttmp834));
AND2X1 AND_tmp836 (.Y(ttmp836),.A(N2779),.B(N2790));
AND2X1 AND_tmp837 (.Y(N7349),.A(N7198),.B(ttmp836));
AND2X1 AND_tmp838 (.Y(ttmp838),.A(N2801),.B(N2812));
AND2X1 AND_tmp839 (.Y(N7357),.A(N7198),.B(ttmp838));
INVX1 NOT1_1886 (.Y(N7363),.A(N7198));
AND2X1 AND_tmp840 (.Y(ttmp840),.A(N1351),.B(N2812));
AND2X1 AND_tmp841 (.Y(N7364),.A(N7190),.B(ttmp840));
INVX1 NOT1_1888 (.Y(N7365),.A(N7190));
NAND2X1 NAND2_1889 (.Y(N7394),.A(N7268),.B(N7184));
NAND2X1 NAND2_1890 (.Y(N7397),.A(N7269),.B(N7186));
NAND2X1 NAND2_1891 (.Y(N7402),.A(N7204),.B(N7300));
INVX1 NOT1_1892 (.Y(N7405),.A(N7209));
NAND2X1 NAND2_1893 (.Y(N7406),.A(N7209),.B(N6884));
INVX1 NOT1_1894 (.Y(N7407),.A(N7212));
NAND2X1 NAND2_1895 (.Y(N7408),.A(N7212),.B(N6888));
NAND2X1 NAND2_1896 (.Y(N7409),.A(N7320),.B(N7216));
NAND2X1 NAND2_1897 (.Y(N7412),.A(N7321),.B(N7218));
INVX1 NOT1_1898 (.Y(N7415),.A(N7219));
NAND2X1 NAND2_1899 (.Y(N7416),.A(N7219),.B(N6904));
INVX1 NOT1_1900 (.Y(N7417),.A(N7222));
NAND2X1 NAND2_1901 (.Y(N7418),.A(N7222),.B(N6908));
INVX1 NOT1_1902 (.Y(N7419),.A(N7225));
NAND2X1 NAND2_1903 (.Y(N7420),.A(N7225),.B(N6913));
NAND2X1 NAND2_1904 (.Y(N7421),.A(N7328),.B(N7229));
INVX1 NOT1_1905 (.Y(N7424),.A(N7245));
INVX1 NOT1_1906 (.Y(N7425),.A(N7242));
INVX1 NOT1_1907 (.Y(N7426),.A(N7239));
INVX1 NOT1_1908 (.Y(N7427),.A(N7236));
INVX1 NOT1_1909 (.Y(N7428),.A(N7263));
INVX1 NOT1_1910 (.Y(N7429),.A(N7260));
INVX1 NOT1_1911 (.Y(N7430),.A(N7257));
INVX1 NOT1_1912 (.Y(N7431),.A(N7250));
INVX1 NOT1_1913 (.Y(N7432),.A(N7250));
AND2X1 AND_tmp842 (.Y(ttmp842),.A(N2653),.B(N2664));
AND2X1 AND_tmp843 (.Y(N7433),.A(N7310),.B(ttmp842));
AND2X1 AND_tmp844 (.Y(ttmp844),.A(N1161),.B(N2664));
AND2X1 AND_tmp845 (.Y(N7434),.A(N7304),.B(ttmp844));
OR2X1 OR_tmp846 (.Y(ttmp846),.A(N3621),.B(N2591));
OR2X1 OR_tmp847 (.Y(ttmp847),.A(N7011),.B(ttmp846));
OR2X1 OR_tmp848 (.Y(N7435),.A(N7338),.B(ttmp847));
AND2X1 AND_tmp849 (.Y(ttmp849),.A(N1185),.B(N2692));
AND2X1 AND_tmp850 (.Y(N7436),.A(N7270),.B(ttmp849));
AND2X1 AND_tmp851 (.Y(ttmp851),.A(N2681),.B(N2692));
AND2X1 AND_tmp852 (.Y(N7437),.A(N7288),.B(ttmp851));
AND2X1 AND_tmp853 (.Y(ttmp853),.A(N1185),.B(N2692));
AND2X1 AND_tmp854 (.Y(N7438),.A(N7276),.B(ttmp853));
AND2X1 AND_tmp855 (.Y(ttmp855),.A(N2681),.B(N2692));
AND2X1 AND_tmp856 (.Y(N7439),.A(N7294),.B(ttmp855));
AND2X1 AND_tmp857 (.Y(ttmp857),.A(N1185),.B(N2692));
AND2X1 AND_tmp858 (.Y(N7440),.A(N7282),.B(ttmp857));
AND2X1 AND_tmp859 (.Y(ttmp859),.A(N2728),.B(N2739));
AND2X1 AND_tmp860 (.Y(N7441),.A(N7310),.B(ttmp859));
AND2X1 AND_tmp861 (.Y(ttmp861),.A(N1223),.B(N2739));
AND2X1 AND_tmp862 (.Y(N7442),.A(N7304),.B(ttmp861));
OR2X1 OR_tmp863 (.Y(ttmp863),.A(N3632),.B(N2600));
OR2X1 OR_tmp864 (.Y(ttmp864),.A(N7012),.B(ttmp863));
OR2X1 OR_tmp865 (.Y(N7443),.A(N7340),.B(ttmp864));
AND2X1 AND_tmp866 (.Y(ttmp866),.A(N1247),.B(N2767));
AND2X1 AND_tmp867 (.Y(N7444),.A(N7270),.B(ttmp866));
AND2X1 AND_tmp868 (.Y(ttmp868),.A(N2756),.B(N2767));
AND2X1 AND_tmp869 (.Y(N7445),.A(N7288),.B(ttmp868));
AND2X1 AND_tmp870 (.Y(ttmp870),.A(N1247),.B(N2767));
AND2X1 AND_tmp871 (.Y(N7446),.A(N7276),.B(ttmp870));
AND2X1 AND_tmp872 (.Y(ttmp872),.A(N2756),.B(N2767));
AND2X1 AND_tmp873 (.Y(N7447),.A(N7294),.B(ttmp872));
AND2X1 AND_tmp874 (.Y(ttmp874),.A(N1247),.B(N2767));
AND2X1 AND_tmp875 (.Y(N7448),.A(N7282),.B(ttmp874));
OR2X1 OR_tmp876 (.Y(ttmp876),.A(N3641),.B(N2605));
OR2X1 OR_tmp877 (.Y(ttmp877),.A(N7013),.B(ttmp876));
OR2X1 OR_tmp878 (.Y(N7449),.A(N7342),.B(ttmp877));
AND2X1 AND_tmp879 (.Y(ttmp879),.A(N3041),.B(N3052));
AND2X1 AND_tmp880 (.Y(N7450),.A(N7310),.B(ttmp879));
AND2X1 AND_tmp881 (.Y(ttmp881),.A(N1697),.B(N3052));
AND2X1 AND_tmp882 (.Y(N7451),.A(N7304),.B(ttmp881));
AND2X1 AND_tmp883 (.Y(ttmp883),.A(N2779),.B(N2790));
AND2X1 AND_tmp884 (.Y(N7452),.A(N7294),.B(ttmp883));
AND2X1 AND_tmp885 (.Y(ttmp885),.A(N1327),.B(N2790));
AND2X1 AND_tmp886 (.Y(N7453),.A(N7282),.B(ttmp885));
AND2X1 AND_tmp887 (.Y(ttmp887),.A(N2779),.B(N2790));
AND2X1 AND_tmp888 (.Y(N7454),.A(N7288),.B(ttmp887));
AND2X1 AND_tmp889 (.Y(ttmp889),.A(N1327),.B(N2790));
AND2X1 AND_tmp890 (.Y(N7455),.A(N7276),.B(ttmp889));
AND2X1 AND_tmp891 (.Y(ttmp891),.A(N1327),.B(N2790));
AND2X1 AND_tmp892 (.Y(N7456),.A(N7270),.B(ttmp891));
AND2X1 AND_tmp893 (.Y(ttmp893),.A(N3075),.B(N3086));
AND2X1 AND_tmp894 (.Y(N7457),.A(N7310),.B(ttmp893));
AND2X1 AND_tmp895 (.Y(ttmp895),.A(N1731),.B(N3086));
AND2X1 AND_tmp896 (.Y(N7458),.A(N7304),.B(ttmp895));
AND2X1 AND_tmp897 (.Y(ttmp897),.A(N2801),.B(N2812));
AND2X1 AND_tmp898 (.Y(N7459),.A(N7294),.B(ttmp897));
AND2X1 AND_tmp899 (.Y(ttmp899),.A(N1351),.B(N2812));
AND2X1 AND_tmp900 (.Y(N7460),.A(N7282),.B(ttmp899));
AND2X1 AND_tmp901 (.Y(ttmp901),.A(N2801),.B(N2812));
AND2X1 AND_tmp902 (.Y(N7461),.A(N7288),.B(ttmp901));
AND2X1 AND_tmp903 (.Y(ttmp903),.A(N1351),.B(N2812));
AND2X1 AND_tmp904 (.Y(N7462),.A(N7276),.B(ttmp903));
AND2X1 AND_tmp905 (.Y(ttmp905),.A(N1351),.B(N2812));
AND2X1 AND_tmp906 (.Y(N7463),.A(N7270),.B(ttmp905));
AND2X1 AND_tmp907 (.Y(ttmp907),.A(N603),.B(N599));
AND2X1 AND_tmp908 (.Y(N7464),.A(N7250),.B(ttmp907));
INVX1 NOT1_1946 (.Y(N7465),.A(N7310));
INVX1 NOT1_1947 (.Y(N7466),.A(N7294));
INVX1 NOT1_1948 (.Y(N7467),.A(N7288));
INVX1 NOT1_1949 (.Y(N7468),.A(N7301));
OR2X1 OR_tmp909 (.Y(ttmp909),.A(N3660),.B(N2626));
OR2X1 OR_tmp910 (.Y(ttmp910),.A(N7016),.B(ttmp909));
OR2X1 OR_tmp911 (.Y(N7469),.A(N7364),.B(ttmp910));
INVX1 NOT1_1951 (.Y(N7470),.A(N7304));
INVX1 NOT1_1952 (.Y(N7471),.A(N7282));
INVX1 NOT1_1953 (.Y(N7472),.A(N7276));
INVX1 NOT1_1954 (.Y(N7473),.A(N7270));
BUFX1 BUFF1_1955 (.Y(N7474),.A(N7394));
BUFX1 BUFF1_1956 (.Y(N7476),.A(N7397));
AND2X1 AND2_1957 (.Y(N7479),.A(N7301),.B(N3068));
AND2X1 AND_tmp912 (.Y(ttmp912),.A(N1793),.B(N3158));
AND2X1 AND_tmp913 (.Y(N7481),.A(N7245),.B(ttmp912));
AND2X1 AND_tmp914 (.Y(ttmp914),.A(N1793),.B(N3158));
AND2X1 AND_tmp915 (.Y(N7482),.A(N7242),.B(ttmp914));
AND2X1 AND_tmp916 (.Y(ttmp916),.A(N1793),.B(N3158));
AND2X1 AND_tmp917 (.Y(N7483),.A(N7239),.B(ttmp916));
AND2X1 AND_tmp918 (.Y(ttmp918),.A(N1793),.B(N3158));
AND2X1 AND_tmp919 (.Y(N7484),.A(N7236),.B(ttmp918));
AND2X1 AND_tmp920 (.Y(ttmp920),.A(N1807),.B(N3180));
AND2X1 AND_tmp921 (.Y(N7485),.A(N7263),.B(ttmp920));
AND2X1 AND_tmp922 (.Y(ttmp922),.A(N1807),.B(N3180));
AND2X1 AND_tmp923 (.Y(N7486),.A(N7260),.B(ttmp922));
AND2X1 AND_tmp924 (.Y(ttmp924),.A(N1807),.B(N3180));
AND2X1 AND_tmp925 (.Y(N7487),.A(N7257),.B(ttmp924));
AND2X1 AND_tmp926 (.Y(ttmp926),.A(N1807),.B(N3180));
AND2X1 AND_tmp927 (.Y(N7488),.A(N7250),.B(ttmp926));
NAND2X1 NAND2_1966 (.Y(N7489),.A(N6979),.B(N7250));
NAND2X1 NAND2_1967 (.Y(N7492),.A(N6516),.B(N7405));
NAND2X1 NAND2_1968 (.Y(N7493),.A(N6526),.B(N7407));
NAND2X1 NAND2_1969 (.Y(N7498),.A(N6592),.B(N7415));
NAND2X1 NAND2_1970 (.Y(N7499),.A(N6599),.B(N7417));
NAND2X1 NAND2_1971 (.Y(N7500),.A(N6609),.B(N7419));
AND2X1 AND_tmp928 (.Y(ttmp928),.A(N7426),.B(N7427));
AND2X1 AND_tmp929 (.Y(ttmp929),.A(N7105),.B(ttmp928));
AND2X1 AND_tmp930 (.Y(ttmp930),.A(N7166),.B(ttmp929));
AND2X1 AND_tmp931 (.Y(ttmp931),.A(N7167),.B(ttmp930));
AND2X1 AND_tmp932 (.Y(ttmp932),.A(N7168),.B(ttmp931));
AND2X1 AND_tmp933 (.Y(ttmp933),.A(N7169),.B(ttmp932));
AND2X1 AND_tmp934 (.Y(ttmp934),.A(N7424),.B(ttmp933));
AND2X1 AND_tmp935 (.Y(N7503),.A(N7425),.B(ttmp934));
AND2X1 AND_tmp936 (.Y(ttmp936),.A(N7430),.B(N7431));
AND2X1 AND_tmp937 (.Y(ttmp937),.A(N6640),.B(ttmp936));
AND2X1 AND_tmp938 (.Y(ttmp938),.A(N7110),.B(ttmp937));
AND2X1 AND_tmp939 (.Y(ttmp939),.A(N7170),.B(ttmp938));
AND2X1 AND_tmp940 (.Y(ttmp940),.A(N7171),.B(ttmp939));
AND2X1 AND_tmp941 (.Y(ttmp941),.A(N7172),.B(ttmp940));
AND2X1 AND_tmp942 (.Y(ttmp942),.A(N7428),.B(ttmp941));
AND2X1 AND_tmp943 (.Y(N7504),.A(N7429),.B(ttmp942));
OR2X1 OR_tmp944 (.Y(ttmp944),.A(N3616),.B(N2585));
OR2X1 OR_tmp945 (.Y(ttmp945),.A(N7433),.B(ttmp944));
OR2X1 OR_tmp946 (.Y(N7505),.A(N7434),.B(ttmp945));
AND2X1 AND2_1975 (.Y(N7506),.A(N7435),.B(N2675));
OR2X1 OR_tmp947 (.Y(ttmp947),.A(N3622),.B(N2592));
OR2X1 OR_tmp948 (.Y(ttmp948),.A(N7339),.B(ttmp947));
OR2X1 OR_tmp949 (.Y(N7507),.A(N7436),.B(ttmp948));
OR2X1 OR_tmp950 (.Y(ttmp950),.A(N3623),.B(N2593));
OR2X1 OR_tmp951 (.Y(ttmp951),.A(N7437),.B(ttmp950));
OR2X1 OR_tmp952 (.Y(N7508),.A(N7438),.B(ttmp951));
OR2X1 OR_tmp953 (.Y(ttmp953),.A(N3624),.B(N2594));
OR2X1 OR_tmp954 (.Y(ttmp954),.A(N7439),.B(ttmp953));
OR2X1 OR_tmp955 (.Y(N7509),.A(N7440),.B(ttmp954));
OR2X1 OR_tmp956 (.Y(ttmp956),.A(N3627),.B(N2595));
OR2X1 OR_tmp957 (.Y(ttmp957),.A(N7441),.B(ttmp956));
OR2X1 OR_tmp958 (.Y(N7510),.A(N7442),.B(ttmp957));
AND2X1 AND2_1980 (.Y(N7511),.A(N7443),.B(N2750));
OR2X1 OR_tmp959 (.Y(ttmp959),.A(N3633),.B(N2601));
OR2X1 OR_tmp960 (.Y(ttmp960),.A(N7341),.B(ttmp959));
OR2X1 OR_tmp961 (.Y(N7512),.A(N7444),.B(ttmp960));
OR2X1 OR_tmp962 (.Y(ttmp962),.A(N3634),.B(N2602));
OR2X1 OR_tmp963 (.Y(ttmp963),.A(N7445),.B(ttmp962));
OR2X1 OR_tmp964 (.Y(N7513),.A(N7446),.B(ttmp963));
OR2X1 OR_tmp965 (.Y(ttmp965),.A(N3635),.B(N2603));
OR2X1 OR_tmp966 (.Y(ttmp966),.A(N7447),.B(ttmp965));
OR2X1 OR_tmp967 (.Y(N7514),.A(N7448),.B(ttmp966));
OR2X1 OR_tmp968 (.Y(ttmp968),.A(N3646),.B(N2610));
OR2X1 OR_tmp969 (.Y(ttmp969),.A(N7450),.B(ttmp968));
OR2X1 OR_tmp970 (.Y(N7515),.A(N7451),.B(ttmp969));
OR2X1 OR_tmp971 (.Y(ttmp971),.A(N3647),.B(N2611));
OR2X1 OR_tmp972 (.Y(ttmp972),.A(N7452),.B(ttmp971));
OR2X1 OR_tmp973 (.Y(N7516),.A(N7453),.B(ttmp972));
OR2X1 OR_tmp974 (.Y(ttmp974),.A(N3648),.B(N2612));
OR2X1 OR_tmp975 (.Y(ttmp975),.A(N7454),.B(ttmp974));
OR2X1 OR_tmp976 (.Y(N7517),.A(N7455),.B(ttmp975));
OR2X1 OR_tmp977 (.Y(ttmp977),.A(N3649),.B(N2613));
OR2X1 OR_tmp978 (.Y(ttmp978),.A(N7349),.B(ttmp977));
OR2X1 OR_tmp979 (.Y(N7518),.A(N7456),.B(ttmp978));
OR2X1 OR_tmp980 (.Y(ttmp980),.A(N3654),.B(N2618));
OR2X1 OR_tmp981 (.Y(ttmp981),.A(N7457),.B(ttmp980));
OR2X1 OR_tmp982 (.Y(N7519),.A(N7458),.B(ttmp981));
OR2X1 OR_tmp983 (.Y(ttmp983),.A(N3655),.B(N2619));
OR2X1 OR_tmp984 (.Y(ttmp984),.A(N7459),.B(ttmp983));
OR2X1 OR_tmp985 (.Y(N7520),.A(N7460),.B(ttmp984));
OR2X1 OR_tmp986 (.Y(ttmp986),.A(N3656),.B(N2620));
OR2X1 OR_tmp987 (.Y(ttmp987),.A(N7461),.B(ttmp986));
OR2X1 OR_tmp988 (.Y(N7521),.A(N7462),.B(ttmp987));
OR2X1 OR_tmp989 (.Y(ttmp989),.A(N3657),.B(N2621));
OR2X1 OR_tmp990 (.Y(ttmp990),.A(N7357),.B(ttmp989));
OR2X1 OR_tmp991 (.Y(N7522),.A(N7463),.B(ttmp990));
OR2X1 OR_tmp992 (.Y(ttmp992),.A(N2624),.B(N7464));
OR2X1 OR_tmp993 (.Y(ttmp993),.A(N4741),.B(ttmp992));
OR2X1 OR_tmp994 (.Y(N7525),.A(N7114),.B(ttmp993));
AND2X1 AND_tmp995 (.Y(ttmp995),.A(N3119),.B(N3130));
AND2X1 AND_tmp996 (.Y(N7526),.A(N7468),.B(ttmp995));
INVX1 NOT1_1994 (.Y(N7527),.A(N7394));
INVX1 NOT1_1995 (.Y(N7528),.A(N7397));
INVX1 NOT1_1996 (.Y(N7529),.A(N7402));
AND2X1 AND2_1997 (.Y(N7530),.A(N7402),.B(N3068));
OR2X1 OR_tmp997 (.Y(ttmp997),.A(N7481),.B(N3801));
OR2X1 OR_tmp998 (.Y(N7531),.A(N4981),.B(ttmp997));
OR2X1 OR_tmp999 (.Y(ttmp999),.A(N7482),.B(N3802));
OR2X1 OR_tmp1000 (.Y(N7537),.A(N4982),.B(ttmp999));
OR2X1 OR_tmp1001 (.Y(ttmp1001),.A(N7483),.B(N3803));
OR2X1 OR_tmp1002 (.Y(N7543),.A(N4983),.B(ttmp1001));
OR2X1 OR_tmp1003 (.Y(ttmp1003),.A(N7484),.B(N3804));
OR2X1 OR_tmp1004 (.Y(N7549),.A(N5165),.B(ttmp1003));
OR2X1 OR_tmp1005 (.Y(ttmp1005),.A(N7485),.B(N3806));
OR2X1 OR_tmp1006 (.Y(N7555),.A(N4985),.B(ttmp1005));
OR2X1 OR_tmp1007 (.Y(ttmp1007),.A(N7486),.B(N3807));
OR2X1 OR_tmp1008 (.Y(N7561),.A(N4986),.B(ttmp1007));
OR2X1 OR_tmp1009 (.Y(ttmp1009),.A(N7487),.B(N3808));
OR2X1 OR_tmp1010 (.Y(N7567),.A(N4547),.B(ttmp1009));
OR2X1 OR_tmp1011 (.Y(ttmp1011),.A(N7488),.B(N3809));
OR2X1 OR_tmp1012 (.Y(N7573),.A(N4987),.B(ttmp1011));
NAND2X1 NAND2_2006 (.Y(N7579),.A(N7492),.B(N7406));
NAND2X1 NAND2_2007 (.Y(N7582),.A(N7493),.B(N7408));
INVX1 NOT1_2008 (.Y(N7585),.A(N7409));
NAND2X1 NAND2_2009 (.Y(N7586),.A(N7409),.B(N6894));
INVX1 NOT1_2010 (.Y(N7587),.A(N7412));
NAND2X1 NAND2_2011 (.Y(N7588),.A(N7412),.B(N6900));
NAND2X1 NAND2_2012 (.Y(N7589),.A(N7498),.B(N7416));
NAND2X1 NAND2_2013 (.Y(N7592),.A(N7499),.B(N7418));
NAND2X1 NAND2_2014 (.Y(N7595),.A(N7500),.B(N7420));
INVX1 NOT1_2015 (.Y(N7598),.A(N7421));
NAND2X1 NAND2_2016 (.Y(N7599),.A(N7421),.B(N6919));
AND2X1 AND2_2017 (.Y(N7600),.A(N7505),.B(N2647));
AND2X1 AND2_2018 (.Y(N7601),.A(N7507),.B(N2675));
AND2X1 AND2_2019 (.Y(N7602),.A(N7508),.B(N2675));
AND2X1 AND2_2020 (.Y(N7603),.A(N7509),.B(N2675));
AND2X1 AND2_2021 (.Y(N7604),.A(N7510),.B(N2722));
AND2X1 AND2_2022 (.Y(N7605),.A(N7512),.B(N2750));
AND2X1 AND2_2023 (.Y(N7606),.A(N7513),.B(N2750));
AND2X1 AND2_2024 (.Y(N7607),.A(N7514),.B(N2750));
AND2X1 AND2_2025 (.Y(N7624),.A(N6979),.B(N7489));
AND2X1 AND2_2026 (.Y(N7625),.A(N7489),.B(N7250));
AND2X1 AND2_2027 (.Y(N7626),.A(N1149),.B(N7525));
AND2X1 AND_tmp1013 (.Y(ttmp1013),.A(N6805),.B(N6930));
AND2X1 AND_tmp1014 (.Y(ttmp1014),.A(N562),.B(ttmp1013));
AND2X1 AND_tmp1015 (.Y(ttmp1015),.A(N7527),.B(ttmp1014));
AND2X1 AND_tmp1016 (.Y(N7631),.A(N7528),.B(ttmp1015));
AND2X1 AND_tmp1017 (.Y(ttmp1017),.A(N3097),.B(N3108));
AND2X1 AND_tmp1018 (.Y(N7636),.A(N7529),.B(ttmp1017));
NAND2X1 NAND2_2030 (.Y(N7657),.A(N6539),.B(N7585));
NAND2X1 NAND2_2031 (.Y(N7658),.A(N6556),.B(N7587));
NAND2X1 NAND2_2032 (.Y(N7665),.A(N6622),.B(N7598));
AND2X1 AND_tmp1019 (.Y(ttmp1019),.A(N2653),.B(N2664));
AND2X1 AND_tmp1020 (.Y(N7666),.A(N7555),.B(ttmp1019));
AND2X1 AND_tmp1021 (.Y(ttmp1021),.A(N1161),.B(N2664));
AND2X1 AND_tmp1022 (.Y(N7667),.A(N7531),.B(ttmp1021));
AND2X1 AND_tmp1023 (.Y(ttmp1023),.A(N2653),.B(N2664));
AND2X1 AND_tmp1024 (.Y(N7668),.A(N7561),.B(ttmp1023));
AND2X1 AND_tmp1025 (.Y(ttmp1025),.A(N1161),.B(N2664));
AND2X1 AND_tmp1026 (.Y(N7669),.A(N7537),.B(ttmp1025));
AND2X1 AND_tmp1027 (.Y(ttmp1027),.A(N2653),.B(N2664));
AND2X1 AND_tmp1028 (.Y(N7670),.A(N7567),.B(ttmp1027));
AND2X1 AND_tmp1029 (.Y(ttmp1029),.A(N1161),.B(N2664));
AND2X1 AND_tmp1030 (.Y(N7671),.A(N7543),.B(ttmp1029));
AND2X1 AND_tmp1031 (.Y(ttmp1031),.A(N2653),.B(N2664));
AND2X1 AND_tmp1032 (.Y(N7672),.A(N7573),.B(ttmp1031));
AND2X1 AND_tmp1033 (.Y(ttmp1033),.A(N1161),.B(N2664));
AND2X1 AND_tmp1034 (.Y(N7673),.A(N7549),.B(ttmp1033));
AND2X1 AND_tmp1035 (.Y(ttmp1035),.A(N2728),.B(N2739));
AND2X1 AND_tmp1036 (.Y(N7674),.A(N7555),.B(ttmp1035));
AND2X1 AND_tmp1037 (.Y(ttmp1037),.A(N1223),.B(N2739));
AND2X1 AND_tmp1038 (.Y(N7675),.A(N7531),.B(ttmp1037));
AND2X1 AND_tmp1039 (.Y(ttmp1039),.A(N2728),.B(N2739));
AND2X1 AND_tmp1040 (.Y(N7676),.A(N7561),.B(ttmp1039));
AND2X1 AND_tmp1041 (.Y(ttmp1041),.A(N1223),.B(N2739));
AND2X1 AND_tmp1042 (.Y(N7677),.A(N7537),.B(ttmp1041));
AND2X1 AND_tmp1043 (.Y(ttmp1043),.A(N2728),.B(N2739));
AND2X1 AND_tmp1044 (.Y(N7678),.A(N7567),.B(ttmp1043));
AND2X1 AND_tmp1045 (.Y(ttmp1045),.A(N1223),.B(N2739));
AND2X1 AND_tmp1046 (.Y(N7679),.A(N7543),.B(ttmp1045));
AND2X1 AND_tmp1047 (.Y(ttmp1047),.A(N2728),.B(N2739));
AND2X1 AND_tmp1048 (.Y(N7680),.A(N7573),.B(ttmp1047));
AND2X1 AND_tmp1049 (.Y(ttmp1049),.A(N1223),.B(N2739));
AND2X1 AND_tmp1050 (.Y(N7681),.A(N7549),.B(ttmp1049));
AND2X1 AND_tmp1051 (.Y(ttmp1051),.A(N3075),.B(N3086));
AND2X1 AND_tmp1052 (.Y(N7682),.A(N7573),.B(ttmp1051));
AND2X1 AND_tmp1053 (.Y(ttmp1053),.A(N1731),.B(N3086));
AND2X1 AND_tmp1054 (.Y(N7683),.A(N7549),.B(ttmp1053));
AND2X1 AND_tmp1055 (.Y(ttmp1055),.A(N3041),.B(N3052));
AND2X1 AND_tmp1056 (.Y(N7684),.A(N7573),.B(ttmp1055));
AND2X1 AND_tmp1057 (.Y(ttmp1057),.A(N1697),.B(N3052));
AND2X1 AND_tmp1058 (.Y(N7685),.A(N7549),.B(ttmp1057));
AND2X1 AND_tmp1059 (.Y(ttmp1059),.A(N3041),.B(N3052));
AND2X1 AND_tmp1060 (.Y(N7686),.A(N7567),.B(ttmp1059));
AND2X1 AND_tmp1061 (.Y(ttmp1061),.A(N1697),.B(N3052));
AND2X1 AND_tmp1062 (.Y(N7687),.A(N7543),.B(ttmp1061));
AND2X1 AND_tmp1063 (.Y(ttmp1063),.A(N3041),.B(N3052));
AND2X1 AND_tmp1064 (.Y(N7688),.A(N7561),.B(ttmp1063));
AND2X1 AND_tmp1065 (.Y(ttmp1065),.A(N1697),.B(N3052));
AND2X1 AND_tmp1066 (.Y(N7689),.A(N7537),.B(ttmp1065));
AND2X1 AND_tmp1067 (.Y(ttmp1067),.A(N3041),.B(N3052));
AND2X1 AND_tmp1068 (.Y(N7690),.A(N7555),.B(ttmp1067));
AND2X1 AND_tmp1069 (.Y(ttmp1069),.A(N1697),.B(N3052));
AND2X1 AND_tmp1070 (.Y(N7691),.A(N7531),.B(ttmp1069));
AND2X1 AND_tmp1071 (.Y(ttmp1071),.A(N3075),.B(N3086));
AND2X1 AND_tmp1072 (.Y(N7692),.A(N7567),.B(ttmp1071));
AND2X1 AND_tmp1073 (.Y(ttmp1073),.A(N1731),.B(N3086));
AND2X1 AND_tmp1074 (.Y(N7693),.A(N7543),.B(ttmp1073));
AND2X1 AND_tmp1075 (.Y(ttmp1075),.A(N3075),.B(N3086));
AND2X1 AND_tmp1076 (.Y(N7694),.A(N7561),.B(ttmp1075));
AND2X1 AND_tmp1077 (.Y(ttmp1077),.A(N1731),.B(N3086));
AND2X1 AND_tmp1078 (.Y(N7695),.A(N7537),.B(ttmp1077));
AND2X1 AND_tmp1079 (.Y(ttmp1079),.A(N3075),.B(N3086));
AND2X1 AND_tmp1080 (.Y(N7696),.A(N7555),.B(ttmp1079));
AND2X1 AND_tmp1081 (.Y(ttmp1081),.A(N1731),.B(N3086));
AND2X1 AND_tmp1082 (.Y(N7697),.A(N7531),.B(ttmp1081));
OR2X1 OR2_2065 (.Y(N7698),.A(N7624),.B(N7625));
INVX1 NOT1_2066 (.Y(N7699),.A(N7573));
INVX1 NOT1_2067 (.Y(N7700),.A(N7567));
INVX1 NOT1_2068 (.Y(N7701),.A(N7561));
INVX1 NOT1_2069 (.Y(N7702),.A(N7555));
AND2X1 AND_tmp1083 (.Y(ttmp1083),.A(N7631),.B(N245));
AND2X1 AND_tmp1084 (.Y(N7703),.A(N1156),.B(ttmp1083));
INVX1 NOT1_2071 (.Y(N7704),.A(N7549));
INVX1 NOT1_2072 (.Y(N7705),.A(N7543));
INVX1 NOT1_2073 (.Y(N7706),.A(N7537));
INVX1 NOT1_2074 (.Y(N7707),.A(N7531));
INVX1 NOT1_2075 (.Y(N7708),.A(N7579));
NAND2X1 NAND2_2076 (.Y(N7709),.A(N7579),.B(N6739));
INVX1 NOT1_2077 (.Y(N7710),.A(N7582));
NAND2X1 NAND2_2078 (.Y(N7711),.A(N7582),.B(N6744));
NAND2X1 NAND2_2079 (.Y(N7712),.A(N7657),.B(N7586));
NAND2X1 NAND2_2080 (.Y(N7715),.A(N7658),.B(N7588));
INVX1 NOT1_2081 (.Y(N7718),.A(N7589));
NAND2X1 NAND2_2082 (.Y(N7719),.A(N7589),.B(N6772));
INVX1 NOT1_2083 (.Y(N7720),.A(N7592));
NAND2X1 NAND2_2084 (.Y(N7721),.A(N7592),.B(N6776));
INVX1 NOT1_2085 (.Y(N7722),.A(N7595));
NAND2X1 NAND2_2086 (.Y(N7723),.A(N7595),.B(N5733));
NAND2X1 NAND2_2087 (.Y(N7724),.A(N7665),.B(N7599));
OR2X1 OR_tmp1085 (.Y(ttmp1085),.A(N3617),.B(N2586));
OR2X1 OR_tmp1086 (.Y(ttmp1086),.A(N7666),.B(ttmp1085));
OR2X1 OR_tmp1087 (.Y(N7727),.A(N7667),.B(ttmp1086));
OR2X1 OR_tmp1088 (.Y(ttmp1088),.A(N3618),.B(N2587));
OR2X1 OR_tmp1089 (.Y(ttmp1089),.A(N7668),.B(ttmp1088));
OR2X1 OR_tmp1090 (.Y(N7728),.A(N7669),.B(ttmp1089));
OR2X1 OR_tmp1091 (.Y(ttmp1091),.A(N3619),.B(N2588));
OR2X1 OR_tmp1092 (.Y(ttmp1092),.A(N7670),.B(ttmp1091));
OR2X1 OR_tmp1093 (.Y(N7729),.A(N7671),.B(ttmp1092));
OR2X1 OR_tmp1094 (.Y(ttmp1094),.A(N3620),.B(N2589));
OR2X1 OR_tmp1095 (.Y(ttmp1095),.A(N7672),.B(ttmp1094));
OR2X1 OR_tmp1096 (.Y(N7730),.A(N7673),.B(ttmp1095));
OR2X1 OR_tmp1097 (.Y(ttmp1097),.A(N3628),.B(N2596));
OR2X1 OR_tmp1098 (.Y(ttmp1098),.A(N7674),.B(ttmp1097));
OR2X1 OR_tmp1099 (.Y(N7731),.A(N7675),.B(ttmp1098));
OR2X1 OR_tmp1100 (.Y(ttmp1100),.A(N3629),.B(N2597));
OR2X1 OR_tmp1101 (.Y(ttmp1101),.A(N7676),.B(ttmp1100));
OR2X1 OR_tmp1102 (.Y(N7732),.A(N7677),.B(ttmp1101));
OR2X1 OR_tmp1103 (.Y(ttmp1103),.A(N3630),.B(N2598));
OR2X1 OR_tmp1104 (.Y(ttmp1104),.A(N7678),.B(ttmp1103));
OR2X1 OR_tmp1105 (.Y(N7733),.A(N7679),.B(ttmp1104));
OR2X1 OR_tmp1106 (.Y(ttmp1106),.A(N3631),.B(N2599));
OR2X1 OR_tmp1107 (.Y(ttmp1107),.A(N7680),.B(ttmp1106));
OR2X1 OR_tmp1108 (.Y(N7734),.A(N7681),.B(ttmp1107));
OR2X1 OR_tmp1109 (.Y(ttmp1109),.A(N3638),.B(N2604));
OR2X1 OR_tmp1110 (.Y(ttmp1110),.A(N7682),.B(ttmp1109));
OR2X1 OR_tmp1111 (.Y(N7735),.A(N7683),.B(ttmp1110));
OR2X1 OR_tmp1112 (.Y(ttmp1112),.A(N3642),.B(N2606));
OR2X1 OR_tmp1113 (.Y(ttmp1113),.A(N7684),.B(ttmp1112));
OR2X1 OR_tmp1114 (.Y(N7736),.A(N7685),.B(ttmp1113));
OR2X1 OR_tmp1115 (.Y(ttmp1115),.A(N3643),.B(N2607));
OR2X1 OR_tmp1116 (.Y(ttmp1116),.A(N7686),.B(ttmp1115));
OR2X1 OR_tmp1117 (.Y(N7737),.A(N7687),.B(ttmp1116));
OR2X1 OR_tmp1118 (.Y(ttmp1118),.A(N3644),.B(N2608));
OR2X1 OR_tmp1119 (.Y(ttmp1119),.A(N7688),.B(ttmp1118));
OR2X1 OR_tmp1120 (.Y(N7738),.A(N7689),.B(ttmp1119));
OR2X1 OR_tmp1121 (.Y(ttmp1121),.A(N3645),.B(N2609));
OR2X1 OR_tmp1122 (.Y(ttmp1122),.A(N7690),.B(ttmp1121));
OR2X1 OR_tmp1123 (.Y(N7739),.A(N7691),.B(ttmp1122));
OR2X1 OR_tmp1124 (.Y(ttmp1124),.A(N3651),.B(N2615));
OR2X1 OR_tmp1125 (.Y(ttmp1125),.A(N7692),.B(ttmp1124));
OR2X1 OR_tmp1126 (.Y(N7740),.A(N7693),.B(ttmp1125));
OR2X1 OR_tmp1127 (.Y(ttmp1127),.A(N3652),.B(N2616));
OR2X1 OR_tmp1128 (.Y(ttmp1128),.A(N7694),.B(ttmp1127));
OR2X1 OR_tmp1129 (.Y(N7741),.A(N7695),.B(ttmp1128));
OR2X1 OR_tmp1130 (.Y(ttmp1130),.A(N3653),.B(N2617));
OR2X1 OR_tmp1131 (.Y(ttmp1131),.A(N7696),.B(ttmp1130));
OR2X1 OR_tmp1132 (.Y(N7742),.A(N7697),.B(ttmp1131));
NAND2X1 NAND2_2104 (.Y(N7743),.A(N6271),.B(N7708));
NAND2X1 NAND2_2105 (.Y(N7744),.A(N6283),.B(N7710));
NAND2X1 NAND2_2106 (.Y(N7749),.A(N6341),.B(N7718));
NAND2X1 NAND2_2107 (.Y(N7750),.A(N6347),.B(N7720));
NAND2X1 NAND2_2108 (.Y(N7751),.A(N5214),.B(N7722));
AND2X1 AND2_2109 (.Y(N7754),.A(N7727),.B(N2647));
AND2X1 AND2_2110 (.Y(N7755),.A(N7728),.B(N2647));
AND2X1 AND2_2111 (.Y(N7756),.A(N7729),.B(N2647));
AND2X1 AND2_2112 (.Y(N7757),.A(N7730),.B(N2647));
AND2X1 AND2_2113 (.Y(N7758),.A(N7731),.B(N2722));
AND2X1 AND2_2114 (.Y(N7759),.A(N7732),.B(N2722));
AND2X1 AND2_2115 (.Y(N7760),.A(N7733),.B(N2722));
AND2X1 AND2_2116 (.Y(N7761),.A(N7734),.B(N2722));
NAND2X1 NAND2_2117 (.Y(N7762),.A(N7743),.B(N7709));
NAND2X1 NAND2_2118 (.Y(N7765),.A(N7744),.B(N7711));
INVX1 NOT1_2119 (.Y(N7768),.A(N7712));
NAND2X1 NAND2_2120 (.Y(N7769),.A(N7712),.B(N6751));
INVX1 NOT1_2121 (.Y(N7770),.A(N7715));
NAND2X1 NAND2_2122 (.Y(N7771),.A(N7715),.B(N6760));
NAND2X1 NAND2_2123 (.Y(N7772),.A(N7749),.B(N7719));
NAND2X1 NAND2_2124 (.Y(N7775),.A(N7750),.B(N7721));
NAND2X1 NAND2_2125 (.Y(N7778),.A(N7751),.B(N7723));
INVX1 NOT1_2126 (.Y(N7781),.A(N7724));
NAND2X1 NAND2_2127 (.Y(N7782),.A(N7724),.B(N5735));
NAND2X1 NAND2_2128 (.Y(N7787),.A(N6295),.B(N7768));
NAND2X1 NAND2_2129 (.Y(N7788),.A(N6313),.B(N7770));
NAND2X1 NAND2_2130 (.Y(N7795),.A(N5220),.B(N7781));
INVX1 NOT1_2131 (.Y(N7796),.A(N7762));
NAND2X1 NAND2_2132 (.Y(N7797),.A(N7762),.B(N6740));
INVX1 NOT1_2133 (.Y(N7798),.A(N7765));
NAND2X1 NAND2_2134 (.Y(N7799),.A(N7765),.B(N6745));
NAND2X1 NAND2_2135 (.Y(N7800),.A(N7787),.B(N7769));
NAND2X1 NAND2_2136 (.Y(N7803),.A(N7788),.B(N7771));
INVX1 NOT1_2137 (.Y(N7806),.A(N7772));
NAND2X1 NAND2_2138 (.Y(N7807),.A(N7772),.B(N6773));
INVX1 NOT1_2139 (.Y(N7808),.A(N7775));
NAND2X1 NAND2_2140 (.Y(N7809),.A(N7775),.B(N6777));
INVX1 NOT1_2141 (.Y(N7810),.A(N7778));
NAND2X1 NAND2_2142 (.Y(N7811),.A(N7778),.B(N6782));
NAND2X1 NAND2_2143 (.Y(N7812),.A(N7795),.B(N7782));
NAND2X1 NAND2_2144 (.Y(N7815),.A(N6274),.B(N7796));
NAND2X1 NAND2_2145 (.Y(N7816),.A(N6286),.B(N7798));
NAND2X1 NAND2_2146 (.Y(N7821),.A(N6344),.B(N7806));
NAND2X1 NAND2_2147 (.Y(N7822),.A(N6350),.B(N7808));
NAND2X1 NAND2_2148 (.Y(N7823),.A(N6353),.B(N7810));
NAND2X1 NAND2_2149 (.Y(N7826),.A(N7815),.B(N7797));
NAND2X1 NAND2_2150 (.Y(N7829),.A(N7816),.B(N7799));
INVX1 NOT1_2151 (.Y(N7832),.A(N7800));
NAND2X1 NAND2_2152 (.Y(N7833),.A(N7800),.B(N6752));
INVX1 NOT1_2153 (.Y(N7834),.A(N7803));
NAND2X1 NAND2_2154 (.Y(N7835),.A(N7803),.B(N6761));
NAND2X1 NAND2_2155 (.Y(N7836),.A(N7821),.B(N7807));
NAND2X1 NAND2_2156 (.Y(N7839),.A(N7822),.B(N7809));
NAND2X1 NAND2_2157 (.Y(N7842),.A(N7823),.B(N7811));
INVX1 NOT1_2158 (.Y(N7845),.A(N7812));
NAND2X1 NAND2_2159 (.Y(N7846),.A(N7812),.B(N6790));
NAND2X1 NAND2_2160 (.Y(N7851),.A(N6298),.B(N7832));
NAND2X1 NAND2_2161 (.Y(N7852),.A(N6316),.B(N7834));
NAND2X1 NAND2_2162 (.Y(N7859),.A(N6364),.B(N7845));
INVX1 NOT1_2163 (.Y(N7860),.A(N7826));
NAND2X1 NAND2_2164 (.Y(N7861),.A(N7826),.B(N6741));
INVX1 NOT1_2165 (.Y(N7862),.A(N7829));
NAND2X1 NAND2_2166 (.Y(N7863),.A(N7829),.B(N6746));
NAND2X1 NAND2_2167 (.Y(N7864),.A(N7851),.B(N7833));
NAND2X1 NAND2_2168 (.Y(N7867),.A(N7852),.B(N7835));
INVX1 NOT1_2169 (.Y(N7870),.A(N7836));
NAND2X1 NAND2_2170 (.Y(N7871),.A(N7836),.B(N5730));
INVX1 NOT1_2171 (.Y(N7872),.A(N7839));
NAND2X1 NAND2_2172 (.Y(N7873),.A(N7839),.B(N5732));
INVX1 NOT1_2173 (.Y(N7874),.A(N7842));
NAND2X1 NAND2_2174 (.Y(N7875),.A(N7842),.B(N6783));
NAND2X1 NAND2_2175 (.Y(N7876),.A(N7859),.B(N7846));
NAND2X1 NAND2_2176 (.Y(N7879),.A(N6277),.B(N7860));
NAND2X1 NAND2_2177 (.Y(N7880),.A(N6289),.B(N7862));
NAND2X1 NAND2_2178 (.Y(N7885),.A(N5199),.B(N7870));
NAND2X1 NAND2_2179 (.Y(N7886),.A(N5208),.B(N7872));
NAND2X1 NAND2_2180 (.Y(N7887),.A(N6356),.B(N7874));
NAND2X1 NAND2_2181 (.Y(N7890),.A(N7879),.B(N7861));
NAND2X1 NAND2_2182 (.Y(N7893),.A(N7880),.B(N7863));
INVX1 NOT1_2183 (.Y(N7896),.A(N7864));
NAND2X1 NAND2_2184 (.Y(N7897),.A(N7864),.B(N6753));
INVX1 NOT1_2185 (.Y(N7898),.A(N7867));
NAND2X1 NAND2_2186 (.Y(N7899),.A(N7867),.B(N6762));
NAND2X1 NAND2_2187 (.Y(N7900),.A(N7885),.B(N7871));
NAND2X1 NAND2_2188 (.Y(N7903),.A(N7886),.B(N7873));
NAND2X1 NAND2_2189 (.Y(N7906),.A(N7887),.B(N7875));
INVX1 NOT1_2190 (.Y(N7909),.A(N7876));
NAND2X1 NAND2_2191 (.Y(N7910),.A(N7876),.B(N6791));
NAND2X1 NAND2_2192 (.Y(N7917),.A(N6301),.B(N7896));
NAND2X1 NAND2_2193 (.Y(N7918),.A(N6319),.B(N7898));
NAND2X1 NAND2_2194 (.Y(N7923),.A(N6367),.B(N7909));
INVX1 NOT1_2195 (.Y(N7924),.A(N7890));
NAND2X1 NAND2_2196 (.Y(N7925),.A(N7890),.B(N6680));
INVX1 NOT1_2197 (.Y(N7926),.A(N7893));
NAND2X1 NAND2_2198 (.Y(N7927),.A(N7893),.B(N6681));
INVX1 NOT1_2199 (.Y(N7928),.A(N7900));
NAND2X1 NAND2_2200 (.Y(N7929),.A(N7900),.B(N5690));
INVX1 NOT1_2201 (.Y(N7930),.A(N7903));
NAND2X1 NAND2_2202 (.Y(N7931),.A(N7903),.B(N5691));
NAND2X1 NAND2_2203 (.Y(N7932),.A(N7917),.B(N7897));
NAND2X1 NAND2_2204 (.Y(N7935),.A(N7918),.B(N7899));
INVX1 NOT1_2205 (.Y(N7938),.A(N7906));
NAND2X1 NAND2_2206 (.Y(N7939),.A(N7906),.B(N6784));
NAND2X1 NAND2_2207 (.Y(N7940),.A(N7923),.B(N7910));
NAND2X1 NAND2_2208 (.Y(N7943),.A(N6280),.B(N7924));
NAND2X1 NAND2_2209 (.Y(N7944),.A(N6292),.B(N7926));
NAND2X1 NAND2_2210 (.Y(N7945),.A(N5202),.B(N7928));
NAND2X1 NAND2_2211 (.Y(N7946),.A(N5211),.B(N7930));
NAND2X1 NAND2_2212 (.Y(N7951),.A(N6359),.B(N7938));
NAND2X1 NAND2_2213 (.Y(N7954),.A(N7943),.B(N7925));
NAND2X1 NAND2_2214 (.Y(N7957),.A(N7944),.B(N7927));
NAND2X1 NAND2_2215 (.Y(N7960),.A(N7945),.B(N7929));
NAND2X1 NAND2_2216 (.Y(N7963),.A(N7946),.B(N7931));
INVX1 NOT1_2217 (.Y(N7966),.A(N7932));
NAND2X1 NAND2_2218 (.Y(N7967),.A(N7932),.B(N6754));
INVX1 NOT1_2219 (.Y(N7968),.A(N7935));
NAND2X1 NAND2_2220 (.Y(N7969),.A(N7935),.B(N6755));
NAND2X1 NAND2_2221 (.Y(N7970),.A(N7951),.B(N7939));
INVX1 NOT1_2222 (.Y(N7973),.A(N7940));
NAND2X1 NAND2_2223 (.Y(N7974),.A(N7940),.B(N6785));
NAND2X1 NAND2_2224 (.Y(N7984),.A(N6304),.B(N7966));
NAND2X1 NAND2_2225 (.Y(N7985),.A(N6322),.B(N7968));
NAND2X1 NAND2_2226 (.Y(N7987),.A(N6370),.B(N7973));
AND2X1 AND_tmp1133 (.Y(ttmp1133),.A(N6831),.B(N1157));
AND2X1 AND_tmp1134 (.Y(N7988),.A(N7957),.B(ttmp1133));
AND2X1 AND_tmp1135 (.Y(ttmp1135),.A(N6415),.B(N1157));
AND2X1 AND_tmp1136 (.Y(N7989),.A(N7954),.B(ttmp1135));
AND2X1 AND_tmp1137 (.Y(ttmp1137),.A(N7041),.B(N566));
AND2X1 AND_tmp1138 (.Y(N7990),.A(N7957),.B(ttmp1137));
AND2X1 AND_tmp1139 (.Y(ttmp1139),.A(N7177),.B(N566));
AND2X1 AND_tmp1140 (.Y(N7991),.A(N7954),.B(ttmp1139));
INVX1 NOT1_2231 (.Y(N7992),.A(N7970));
NAND2X1 NAND2_2232 (.Y(N7993),.A(N7970),.B(N6448));
AND2X1 AND_tmp1141 (.Y(ttmp1141),.A(N6857),.B(N1219));
AND2X1 AND_tmp1142 (.Y(N7994),.A(N7963),.B(ttmp1141));
AND2X1 AND_tmp1143 (.Y(ttmp1143),.A(N6441),.B(N1219));
AND2X1 AND_tmp1144 (.Y(N7995),.A(N7960),.B(ttmp1143));
AND2X1 AND_tmp1145 (.Y(ttmp1145),.A(N7065),.B(N583));
AND2X1 AND_tmp1146 (.Y(N7996),.A(N7963),.B(ttmp1145));
AND2X1 AND_tmp1147 (.Y(ttmp1147),.A(N7182),.B(N583));
AND2X1 AND_tmp1148 (.Y(N7997),.A(N7960),.B(ttmp1147));
NAND2X1 NAND2_2237 (.Y(N7998),.A(N7984),.B(N7967));
NAND2X1 NAND2_2238 (.Y(N8001),.A(N7985),.B(N7969));
NAND2X1 NAND2_2239 (.Y(N8004),.A(N7987),.B(N7974));
NAND2X1 NAND2_2240 (.Y(N8009),.A(N6051),.B(N7992));
OR2X1 OR_tmp1149 (.Y(ttmp1149),.A(N7990),.B(N7991));
OR2X1 OR_tmp1150 (.Y(ttmp1150),.A(N7988),.B(ttmp1149));
OR2X1 OR_tmp1151 (.Y(N8013),.A(N7989),.B(ttmp1150));
OR2X1 OR_tmp1152 (.Y(ttmp1152),.A(N7996),.B(N7997));
OR2X1 OR_tmp1153 (.Y(ttmp1153),.A(N7994),.B(ttmp1152));
OR2X1 OR_tmp1154 (.Y(N8017),.A(N7995),.B(ttmp1153));
INVX1 NOT1_2243 (.Y(N8020),.A(N7998));
NAND2X1 NAND2_2244 (.Y(N8021),.A(N7998),.B(N6682));
INVX1 NOT1_2245 (.Y(N8022),.A(N8001));
NAND2X1 NAND2_2246 (.Y(N8023),.A(N8001),.B(N6683));
NAND2X1 NAND2_2247 (.Y(N8025),.A(N8009),.B(N7993));
INVX1 NOT1_2248 (.Y(N8026),.A(N8004));
NAND2X1 NAND2_2249 (.Y(N8027),.A(N8004),.B(N6449));
NAND2X1 NAND2_2250 (.Y(N8031),.A(N6307),.B(N8020));
NAND2X1 NAND2_2251 (.Y(N8032),.A(N6310),.B(N8022));
INVX1 NOT1_2252 (.Y(N8033),.A(N8013));
NAND2X1 NAND2_2253 (.Y(N8034),.A(N6054),.B(N8026));
AND2X1 AND2_2254 (.Y(N8035),.A(N583),.B(N8025));
INVX1 NOT1_2255 (.Y(N8036),.A(N8017));
NAND2X1 NAND2_2256 (.Y(N8037),.A(N8031),.B(N8021));
NAND2X1 NAND2_2257 (.Y(N8038),.A(N8032),.B(N8023));
NAND2X1 NAND2_2258 (.Y(N8039),.A(N8034),.B(N8027));
INVX1 NOT1_2259 (.Y(N8040),.A(N8038));
AND2X1 AND2_2260 (.Y(N8041),.A(N566),.B(N8037));
INVX1 NOT1_2261 (.Y(N8042),.A(N8039));
AND2X1 AND2_2262 (.Y(N8043),.A(N8040),.B(N1157));
AND2X1 AND2_2263 (.Y(N8044),.A(N8042),.B(N1219));
OR2X1 OR2_2264 (.Y(N8045),.A(N8043),.B(N8041));
OR2X1 OR2_2265 (.Y(N8048),.A(N8044),.B(N8035));
NAND2X1 NAND2_2266 (.Y(N8055),.A(N8045),.B(N8033));
INVX1 NOT1_2267 (.Y(N8056),.A(N8045));
NAND2X1 NAND2_2268 (.Y(N8057),.A(N8048),.B(N8036));
INVX1 NOT1_2269 (.Y(N8058),.A(N8048));
NAND2X1 NAND2_2270 (.Y(N8059),.A(N8013),.B(N8056));
NAND2X1 NAND2_2271 (.Y(N8060),.A(N8017),.B(N8058));
NAND2X1 NAND2_2272 (.Y(N8061),.A(N8055),.B(N8059));
NAND2X1 NAND2_2273 (.Y(N8064),.A(N8057),.B(N8060));
AND2X1 AND_tmp1155 (.Y(ttmp1155),.A(N1777),.B(N3130));
AND2X1 AND_tmp1156 (.Y(N8071),.A(N8064),.B(ttmp1155));
AND2X1 AND_tmp1157 (.Y(ttmp1157),.A(N1761),.B(N3108));
AND2X1 AND_tmp1158 (.Y(N8072),.A(N8061),.B(ttmp1157));
INVX1 NOT1_2276 (.Y(N8073),.A(N8061));
INVX1 NOT1_2277 (.Y(N8074),.A(N8064));
OR2X1 OR_tmp1159 (.Y(ttmp1159),.A(N3659),.B(N2625));
OR2X1 OR_tmp1160 (.Y(ttmp1160),.A(N7526),.B(ttmp1159));
OR2X1 OR_tmp1161 (.Y(N8075),.A(N8071),.B(ttmp1160));
OR2X1 OR_tmp1162 (.Y(ttmp1162),.A(N3661),.B(N2627));
OR2X1 OR_tmp1163 (.Y(ttmp1163),.A(N7636),.B(ttmp1162));
OR2X1 OR_tmp1164 (.Y(N8076),.A(N8072),.B(ttmp1163));
AND2X1 AND2_2280 (.Y(N8077),.A(N8073),.B(N1727));
AND2X1 AND2_2281 (.Y(N8078),.A(N8074),.B(N1727));
OR2X1 OR2_2282 (.Y(N8079),.A(N7530),.B(N8077));
OR2X1 OR2_2283 (.Y(N8082),.A(N7479),.B(N8078));
AND2X1 AND2_2284 (.Y(N8089),.A(N8079),.B(N3063));
AND2X1 AND2_2285 (.Y(N8090),.A(N8082),.B(N3063));
AND2X1 AND2_2286 (.Y(N8091),.A(N8079),.B(N3063));
AND2X1 AND2_2287 (.Y(N8092),.A(N8082),.B(N3063));
OR2X1 OR2_2288 (.Y(N8093),.A(N8089),.B(N3071));
OR2X1 OR2_2289 (.Y(N8096),.A(N8090),.B(N3072));
OR2X1 OR2_2290 (.Y(N8099),.A(N8091),.B(N3073));
OR2X1 OR2_2291 (.Y(N8102),.A(N8092),.B(N3074));
AND2X1 AND_tmp1165 (.Y(ttmp1165),.A(N2779),.B(N2790));
AND2X1 AND_tmp1166 (.Y(N8113),.A(N8102),.B(ttmp1165));
AND2X1 AND_tmp1167 (.Y(ttmp1167),.A(N1327),.B(N2790));
AND2X1 AND_tmp1168 (.Y(N8114),.A(N8099),.B(ttmp1167));
AND2X1 AND_tmp1169 (.Y(ttmp1169),.A(N2801),.B(N2812));
AND2X1 AND_tmp1170 (.Y(N8115),.A(N8102),.B(ttmp1169));
AND2X1 AND_tmp1171 (.Y(ttmp1171),.A(N1351),.B(N2812));
AND2X1 AND_tmp1172 (.Y(N8116),.A(N8099),.B(ttmp1171));
AND2X1 AND_tmp1173 (.Y(ttmp1173),.A(N2681),.B(N2692));
AND2X1 AND_tmp1174 (.Y(N8117),.A(N8096),.B(ttmp1173));
AND2X1 AND_tmp1175 (.Y(ttmp1175),.A(N1185),.B(N2692));
AND2X1 AND_tmp1176 (.Y(N8118),.A(N8093),.B(ttmp1175));
AND2X1 AND_tmp1177 (.Y(ttmp1177),.A(N2756),.B(N2767));
AND2X1 AND_tmp1178 (.Y(N8119),.A(N8096),.B(ttmp1177));
AND2X1 AND_tmp1179 (.Y(ttmp1179),.A(N1247),.B(N2767));
AND2X1 AND_tmp1180 (.Y(N8120),.A(N8093),.B(ttmp1179));
OR2X1 OR_tmp1181 (.Y(ttmp1181),.A(N3662),.B(N2703));
OR2X1 OR_tmp1182 (.Y(ttmp1182),.A(N8117),.B(ttmp1181));
OR2X1 OR_tmp1183 (.Y(N8121),.A(N8118),.B(ttmp1182));
OR2X1 OR_tmp1184 (.Y(ttmp1184),.A(N3663),.B(N2778));
OR2X1 OR_tmp1185 (.Y(ttmp1185),.A(N8119),.B(ttmp1184));
OR2X1 OR_tmp1186 (.Y(N8122),.A(N8120),.B(ttmp1185));
OR2X1 OR_tmp1187 (.Y(ttmp1187),.A(N3650),.B(N2614));
OR2X1 OR_tmp1188 (.Y(ttmp1188),.A(N8113),.B(ttmp1187));
OR2X1 OR_tmp1189 (.Y(N8123),.A(N8114),.B(ttmp1188));
OR2X1 OR_tmp1190 (.Y(ttmp1190),.A(N3658),.B(N2622));
OR2X1 OR_tmp1191 (.Y(ttmp1191),.A(N8115),.B(ttmp1190));
OR2X1 OR_tmp1192 (.Y(N8124),.A(N8116),.B(ttmp1191));
AND2X1 AND2_2304 (.Y(N8125),.A(N8121),.B(N2675));
AND2X1 AND2_2305 (.Y(N8126),.A(N8122),.B(N2750));
INVX1 NOT1_2306 (.Y(N8127),.A(N8125));
INVX1 NOT1_2307 (.Y(N8128),.A(N8126));
XNOR2X1 compare_0 (.Y(compare0),.A(keyinput0),.B(N1));
XNOR2X1 compare_1 (.Y(compare1),.A(keyinput1),.B(N4));
XNOR2X1 compare_2 (.Y(compare2),.A(keyinput2),.B(N11));
XNOR2X1 compare_3 (.Y(compare3),.A(keyinput3),.B(N14));
XNOR2X1 compare_4 (.Y(compare4),.A(keyinput4),.B(N17));
XNOR2X1 compare_5 (.Y(compare5),.A(keyinput5),.B(N20));
XNOR2X1 compare_6 (.Y(compare6),.A(keyinput6),.B(N23));
XNOR2X1 compare_7 (.Y(compare7),.A(keyinput7),.B(N24));
XNOR2X1 compare_8 (.Y(compare8),.A(keyinput8),.B(N25));
XNOR2X1 compare_9 (.Y(compare9),.A(keyinput9),.B(N26));
XNOR2X1 compare_10 (.Y(compare10),.A(keyinput10),.B(N27));
XNOR2X1 compare_11 (.Y(compare11),.A(keyinput11),.B(N31));
AND2X1 andgate_0 (.Y(andgate0),.A(compare0),.B(compare1));
AND2X1 andgate_1 (.Y(andgate1),.A(compare2),.B(compare3));
AND2X1 andgate_2 (.Y(andgate2),.A(compare4),.B(compare5));
AND2X1 andgate_3 (.Y(andgate3),.A(compare6),.B(compare7));
AND2X1 andgate_4 (.Y(andgate4),.A(compare8),.B(compare9));
AND2X1 andgate_5 (.Y(andgate5),.A(compare10),.B(compare11));
AND2X1 andgate_6 (.Y(andgate6),.A(andgate0),.B(andgate1));
AND2X1 andgate_7 (.Y(andgate7),.A(andgate2),.B(andgate3));
AND2X1 andgate_8 (.Y(andgate8),.A(andgate4),.B(andgate5));
AND2X1 andgate_9 (.Y(andgate9),.A(andgate6),.B(andgate7));
AND2X1 andgate_10 (.Y(andgate10),.A(andgate8),.B(andgate9));
OR2X1 orgate_0 (.Y(orgate0),.A(keyinput0),.B(keyinput1));
OR2X1 orgate_1 (.Y(orgate1),.A(keyinput2),.B(keyinput3));
OR2X1 orgate_2 (.Y(orgate2),.A(keyinput4),.B(keyinput5));
OR2X1 orgate_3 (.Y(orgate3),.A(keyinput6),.B(keyinput7));
OR2X1 orgate_4 (.Y(orgate4),.A(keyinput8),.B(keyinput9));
OR2X1 orgate_5 (.Y(orgate5),.A(keyinput10),.B(keyinput11));
OR2X1 orgate_6 (.Y(orgate6),.A(orgate0),.B(orgate1));
OR2X1 orgate_7 (.Y(orgate7),.A(orgate2),.B(orgate3));
OR2X1 orgate_8 (.Y(orgate8),.A(orgate4),.B(orgate5));
OR2X1 orgate_9 (.Y(orgate9),.A(orgate6),.B(orgate7));
OR2X1 orgate_10 (.Y(orgate10),.A(orgate8),.B(orgate9));
AND2X1 andgate_11 (.Y(andgate11),.A(orgate10),.B(andgate10));
XOR2X1 XOR_out0 (.Y(N709),.A(N709_sar),.B(andgate11));
endmodule