module c7552 (N1,N5,N9,N12,N15,N18,N23,N26,N29,N32,N35,N38,N41,N44,N47,N50,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N69,N70,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N94,N97,N100,N103,N106,N109,N110,N111,N112,N113,N114,N115,N118,N121,N124,N127,N130,N133,N134,N135,N138,N141,N144,N147,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N242,N245,N248,N251,N254,N257,N260,N263,N267,N271,N274,N277,N280,N283,N286,N289,N293,N296,N299,N303,N307,N310,N313,N316,N319,N322,N325,N328,N331,N334,N337,N340,N343,N346,N349,N352,N355,N358,N361,N364,N367,N382,N241_I,N387,N388,N478,N482,N484,N486,N489,N492,N501,N505,N507,N509,N511,N513,N515,N517,N519,N535,N537,N539,N541,N543,N545,N547,N549,N551,N553,N556,N559,N561,N563,N565,N567,N569,N571,N573,N582,N643,N707,N813,N881,N882,N883,N884,N885,N889,N945,N1110,N1111,N1112,N1113,N1114,N1489,N1490,N1781,N10025,N10101,N10102,N10103,N10104,N10109,N10110,N10111,N10112,N10350,N10351,N10352,N10353,N10574,N10575,N10576,N10628,N10632,N10641,N10704,N10706,N10711,N10712,N10713,N10714,N10715,N10716,N10717,N10718,N10729,N10759,N10760,N10761,N10762,N10763,N10827,N10837,N10838,N10839,N10840,N10868,N10869,N10870,N10871,N10905,N10906,N10907,N10908,N11333,N11334,N11340,N11342,N241_O);
input N1,N5,N9,N12,N15,N18,N23,N26,N29,N32,N35,N38,N41,N44,N47,N50,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N69,N70,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N94,N97,N100,N103,N106,N109,N110,N111,N112,N113,N114,N115,N118,N121,N124,N127,N130,N133,N134,N135,N138,N141,N144,N147,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N242,N245,N248,N251,N254,N257,N260,N263,N267,N271,N274,N277,N280,N283,N286,N289,N293,N296,N299,N303,N307,N310,N313,N316,N319,N322,N325,N328,N331,N334,N337,N340,N343,N346,N349,N352,N355,N358,N361,N364,N367,N382,N241_I;
output N387,N388,N478,N482,N484,N486,N489,N492,N501,N505,N507,N509,N511,N513,N515,N517,N519,N535,N537,N539,N541,N543,N545,N547,N549,N551,N553,N556,N559,N561,N563,N565,N567,N569,N571,N573,N582,N643,N707,N813,N881,N882,N883,N884,N885,N889,N945,N1110,N1111,N1112,N1113,N1114,N1489,N1490,N1781,N10025,N10101,N10102,N10103,N10104,N10109,N10110,N10111,N10112,N10350,N10351,N10352,N10353,N10574,N10575,N10576,N10628,N10632,N10641,N10704,N10706,N10711,N10712,N10713,N10714,N10715,N10716,N10717,N10718,N10729,N10759,N10760,N10761,N10762,N10763,N10827,N10837,N10838,N10839,N10840,N10868,N10869,N10870,N10871,N10905,N10906,N10907,N10908,N11333,N11334,N11340,N11342,N241_O;
wire N467,N469,N494,N528,N575,N578,N585,N590,N593,N596,N599,N604,N609,N614,N625,N628,N632,N636,N641,N642,N644,N651,N657,N660,N666,N672,N673,N674,N676,N682,N688,N689,N695,N700,N705,N706,N708,N715,N721,N727,N733,N734,N742,N748,N749,N750,N758,N759,N762,N768,N774,N780,N786,N794,N800,N806,N812,N814,N821,N827,N833,N839,N845,N853,N859,N865,N871,N886,N887,N957,N1028,N1029,N1109,N1115,N1116,N1119,N1125,N1132,N1136,N1141,N1147,N1154,N1160,N1167,N1174,N1175,N1182,N1189,N1194,N1199,N1206,N1211,N1218,N1222,N1227,N1233,N1240,N1244,N1249,N1256,N1263,N1270,N1277,N1284,N1287,N1290,N1293,N1296,N1299,N1302,N1305,N1308,N1311,N1314,N1317,N1320,N1323,N1326,N1329,N1332,N1335,N1338,N1341,N1344,N1347,N1350,N1353,N1356,N1359,N1362,N1365,N1368,N1371,N1374,N1377,N1380,N1383,N1386,N1389,N1392,N1395,N1398,N1401,N1404,N1407,N1410,N1413,N1416,N1419,N1422,N1425,N1428,N1431,N1434,N1437,N1440,N1443,N1446,N1449,N1452,N1455,N1458,N1461,N1464,N1467,N1470,N1473,N1476,N1479,N1482,N1485,N1537,N1551,N1649,N1703,N1708,N1713,N1721,N1758,N1782,N1783,N1789,N1793,N1794,N1795,N1796,N1797,N1798,N1799,N1805,N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,N1819,N1820,N1821,N1822,N1828,N1829,N1830,N1832,N1833,N1834,N1835,N1839,N1840,N1841,N1842,N1843,N1845,N1851,N1857,N1858,N1859,N1860,N1861,N1862,N1863,N1864,N1865,N1866,N1867,N1868,N1869,N1870,N1871,N1872,N1873,N1874,N1875,N1876,N1877,N1878,N1879,N1880,N1881,N1882,N1883,N1884,N1885,N1892,N1899,N1906,N1913,N1919,N1926,N1927,N1928,N1929,N1930,N1931,N1932,N1933,N1934,N1935,N1936,N1937,N1938,N1939,N1940,N1941,N1942,N1943,N1944,N1945,N1946,N1947,N1953,N1957,N1958,N1959,N1960,N1961,N1962,N1963,N1965,N1966,N1967,N1968,N1969,N1970,N1971,N1972,N1973,N1974,N1975,N1976,N1977,N1983,N1989,N1990,N1991,N1992,N1993,N1994,N1995,N1996,N1997,N2003,N2010,N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,N2019,N2020,N2021,N2022,N2023,N2024,N2031,N2038,N2045,N2052,N2058,N2064,N2065,N2066,N2067,N2068,N2069,N2070,N2071,N2072,N2073,N2074,N2081,N2086,N2107,N2108,N2110,N2111,N2112,N2113,N2114,N2115,N2117,N2171,N2172,N2230,N2231,N2235,N2239,N2240,N2241,N2242,N2243,N2244,N2245,N2246,N2247,N2248,N2249,N2250,N2251,N2252,N2253,N2254,N2255,N2256,N2257,N2267,N2268,N2269,N2274,N2275,N2277,N2278,N2279,N2280,N2281,N2282,N2283,N2284,N2285,N2286,N2287,N2293,N2299,N2300,N2301,N2302,N2303,N2304,N2305,N2306,N2307,N2308,N2309,N2315,N2321,N2322,N2323,N2324,N2325,N2326,N2327,N2328,N2329,N2330,N2331,N2337,N2338,N2339,N2340,N2341,N2342,N2343,N2344,N2345,N2346,N2347,N2348,N2349,N2350,N2351,N2352,N2353,N2354,N2355,N2356,N2357,N2358,N2359,N2360,N2361,N2362,N2363,N2364,N2365,N2366,N2367,N2368,N2374,N2375,N2376,N2377,N2378,N2379,N2380,N2381,N2382,N2383,N2384,N2390,N2396,N2397,N2398,N2399,N2400,N2401,N2402,N2403,N2404,N2405,N2406,N2412,N2418,N2419,N2420,N2421,N2422,N2423,N2424,N2425,N2426,N2427,N2428,N2429,N2430,N2431,N2432,N2433,N2434,N2435,N2436,N2437,N2441,N2442,N2446,N2450,N2454,N2458,N2462,N2466,N2470,N2474,N2478,N2482,N2488,N2496,N2502,N2508,N2523,N2533,N2537,N2538,N2542,N2546,N2550,N2554,N2561,N2567,N2573,N2604,N2607,N2611,N2615,N2619,N2626,N2632,N2638,N2644,N2650,N2653,N2654,N2658,N2662,N2666,N2670,N2674,N2680,N2688,N2692,N2696,N2700,N2704,N2728,N2729,N2733,N2737,N2741,N2745,N2749,N2753,N2757,N2761,N2765,N2766,N2769,N2772,N2775,N2778,N2781,N2784,N2787,N2790,N2793,N2796,N2866,N2867,N2868,N2869,N2878,N2913,N2914,N2915,N2916,N2917,N2918,N2919,N2920,N2921,N2922,N2923,N2924,N2925,N2926,N2927,N2928,N2929,N2930,N2931,N2932,N2933,N2934,N2935,N2936,N2937,N2988,N3005,N3006,N3007,N3008,N3009,N3020,N3021,N3022,N3023,N3024,N3025,N3026,N3027,N3028,N3029,N3032,N3033,N3034,N3035,N3036,N3037,N3038,N3039,N3040,N3041,N3061,N3064,N3067,N3070,N3073,N3080,N3096,N3097,N3101,N3107,N3114,N3122,N3126,N3130,N3131,N3134,N3135,N3136,N3137,N3140,N3144,N3149,N3155,N3159,N3167,N3168,N3169,N3173,N3178,N3184,N3185,N3189,N3195,N3202,N3210,N3211,N3215,N3221,N3228,N3229,N3232,N3236,N3241,N3247,N3251,N3255,N3259,N3263,N3267,N3273,N3281,N3287,N3293,N3299,N3303,N3307,N3311,N3315,N3322,N3328,N3334,N3340,N3343,N3349,N3355,N3361,N3362,N3363,N3364,N3365,N3366,N3367,N3368,N3369,N3370,N3371,N3372,N3373,N3374,N3375,N3379,N3380,N3381,N3384,N3390,N3398,N3404,N3410,N3416,N3420,N3424,N3428,N3432,N3436,N3440,N3444,N3448,N3452,N3453,N3454,N3458,N3462,N3466,N3470,N3474,N3478,N3482,N3486,N3487,N3490,N3493,N3496,N3499,N3502,N3507,N3510,N3515,N3518,N3521,N3524,N3527,N3530,N3535,N3539,N3542,N3545,N3548,N3551,N3552,N3553,N3557,N3560,N3563,N3566,N3569,N3570,N3571,N3574,N3577,N3580,N3583,N3586,N3589,N3592,N3595,N3598,N3601,N3604,N3607,N3610,N3613,N3616,N3619,N3622,N3625,N3628,N3631,N3634,N3637,N3640,N3643,N3646,N3649,N3652,N3655,N3658,N3661,N3664,N3667,N3670,N3673,N3676,N3679,N3682,N3685,N3688,N3691,N3694,N3697,N3700,N3703,N3706,N3709,N3712,N3715,N3718,N3721,N3724,N3727,N3730,N3733,N3736,N3739,N3742,N3745,N3748,N3751,N3754,N3757,N3760,N3763,N3766,N3769,N3772,N3775,N3778,N3781,N3782,N3783,N3786,N3789,N3792,N3795,N3798,N3801,N3804,N3807,N3810,N3813,N3816,N3819,N3822,N3825,N3828,N3831,N3834,N3837,N3840,N3843,N3846,N3849,N3852,N3855,N3858,N3861,N3864,N3867,N3870,N3873,N3876,N3879,N3882,N3885,N3888,N3891,N3953,N3954,N3955,N3956,N3958,N3964,N4193,N4303,N4308,N4313,N4326,N4327,N4333,N4334,N4411,N4412,N4463,N4464,N4465,N4466,N4467,N4468,N4469,N4470,N4471,N4472,N4473,N4474,N4475,N4476,N4477,N4478,N4479,N4480,N4481,N4482,N4483,N4484,N4485,N4486,N4487,N4488,N4489,N4490,N4491,N4492,N4493,N4494,N4495,N4496,N4497,N4498,N4499,N4500,N4501,N4502,N4503,N4504,N4505,N4506,N4507,N4508,N4509,N4510,N4511,N4512,N4513,N4514,N4515,N4516,N4517,N4518,N4519,N4520,N4521,N4522,N4523,N4524,N4525,N4526,N4527,N4528,N4529,N4530,N4531,N4532,N4533,N4534,N4535,N4536,N4537,N4538,N4539,N4540,N4541,N4542,N4543,N4544,N4545,N4549,N4555,N4562,N4563,N4566,N4570,N4575,N4576,N4577,N4581,N4586,N4592,N4593,N4597,N4603,N4610,N4611,N4612,N4613,N4614,N4615,N4616,N4617,N4618,N4619,N4620,N4621,N4622,N4623,N4624,N4625,N4626,N4627,N4628,N4629,N4630,N4631,N4632,N4633,N4634,N4635,N4636,N4637,N4638,N4639,N4640,N4641,N4642,N4643,N4644,N4645,N4646,N4647,N4648,N4649,N4650,N4651,N4652,N4653,N4656,N4657,N4661,N4667,N4674,N4675,N4678,N4682,N4687,N4693,N4694,N4695,N4696,N4697,N4698,N4699,N4700,N4701,N4702,N4706,N4711,N4717,N4718,N4722,N4728,N4735,N4743,N4744,N4745,N4746,N4747,N4748,N4749,N4750,N4751,N4752,N4753,N4754,N4755,N4756,N4757,N4758,N4759,N4760,N4761,N4762,N4763,N4764,N4765,N4766,N4767,N4768,N4769,N4775,N4776,N4777,N4778,N4779,N4780,N4781,N4782,N4783,N4784,N4789,N4790,N4793,N4794,N4795,N4796,N4799,N4800,N4801,N4802,N4803,N4806,N4809,N4810,N4813,N4814,N4817,N4820,N4823,N4826,N4829,N4832,N4835,N4838,N4841,N4844,N4847,N4850,N4853,N4856,N4859,N4862,N4865,N4868,N4871,N4874,N4877,N4880,N4883,N4886,N4889,N4892,N4895,N4898,N4901,N4904,N4907,N4910,N4913,N4916,N4919,N4922,N4925,N4928,N4931,N4934,N4937,N4940,N4943,N4946,N4949,N4952,N4955,N4958,N4961,N4964,N4967,N4970,N4973,N4976,N4979,N4982,N4985,N4988,N4991,N4994,N4997,N5000,N5003,N5006,N5009,N5012,N5015,N5018,N5021,N5024,N5027,N5030,N5033,N5036,N5039,N5042,N5045,N5046,N5047,N5048,N5049,N5052,N5055,N5058,N5061,N5064,N5065,N5066,N5067,N5068,N5071,N5074,N5077,N5080,N5083,N5086,N5089,N5092,N5095,N5098,N5101,N5104,N5107,N5110,N5111,N5112,N5113,N5114,N5117,N5120,N5123,N5126,N5129,N5132,N5135,N5138,N5141,N5144,N5147,N5150,N5153,N5156,N5159,N5162,N5165,N5166,N5167,N5168,N5169,N5170,N5171,N5172,N5173,N5174,N5175,N5176,N5177,N5178,N5179,N5180,N5181,N5182,N5183,N5184,N5185,N5186,N5187,N5188,N5189,N5190,N5191,N5192,N5193,N5196,N5197,N5198,N5199,N5200,N5201,N5202,N5203,N5204,N5205,N5206,N5207,N5208,N5209,N5210,N5211,N5212,N5213,N5283,N5284,N5285,N5286,N5287,N5288,N5289,N5290,N5291,N5292,N5293,N5294,N5295,N5296,N5297,N5298,N5299,N5300,N5314,N5315,N5316,N5317,N5318,N5319,N5320,N5321,N5322,N5323,N5324,N5363,N5364,N5365,N5366,N5367,N5425,N5426,N5427,N5429,N5430,N5431,N5432,N5433,N5451,N5452,N5453,N5454,N5455,N5456,N5457,N5469,N5474,N5475,N5476,N5477,N5571,N5572,N5573,N5574,N5584,N5585,N5586,N5587,N5602,N5603,N5604,N5605,N5631,N5632,N5640,N5654,N5670,N5683,N5690,N5697,N5707,N5718,N5728,N5735,N5736,N5740,N5744,N5747,N5751,N5755,N5758,N5762,N5766,N5769,N5770,N5771,N5778,N5789,N5799,N5807,N5821,N5837,N5850,N5856,N5863,N5870,N5881,N5892,N5898,N5905,N5915,N5926,N5936,N5943,N5944,N5945,N5946,N5947,N5948,N5949,N5950,N5951,N5952,N5953,N5954,N5955,N5956,N5957,N5958,N5959,N5960,N5966,N5967,N5968,N5969,N5970,N5971,N5972,N5973,N5974,N5975,N5976,N5977,N5978,N5979,N5980,N5981,N5989,N5990,N5991,N5996,N6000,N6003,N6009,N6014,N6018,N6021,N6022,N6023,N6024,N6025,N6026,N6027,N6028,N6029,N6030,N6031,N6032,N6033,N6034,N6035,N6036,N6037,N6038,N6039,N6040,N6041,N6047,N6052,N6056,N6059,N6060,N6061,N6062,N6063,N6064,N6065,N6066,N6067,N6068,N6069,N6070,N6071,N6072,N6073,N6074,N6075,N6076,N6077,N6078,N6079,N6083,N6087,N6090,N6091,N6092,N6093,N6094,N6095,N6096,N6097,N6098,N6099,N6100,N6101,N6102,N6103,N6104,N6105,N6106,N6107,N6108,N6109,N6110,N6111,N6112,N6113,N6114,N6115,N6116,N6117,N6118,N6119,N6120,N6121,N6122,N6123,N6124,N6125,N6126,N6127,N6131,N6135,N6136,N6137,N6141,N6145,N6148,N6149,N6150,N6151,N6152,N6153,N6154,N6155,N6156,N6157,N6158,N6159,N6160,N6161,N6162,N6163,N6164,N6165,N6166,N6170,N6174,N6177,N6181,N6182,N6183,N6184,N6185,N6186,N6187,N6188,N6189,N6190,N6191,N6192,N6193,N6194,N6195,N6196,N6199,N6202,N6203,N6204,N6207,N6210,N6213,N6214,N6217,N6220,N6223,N6224,N6225,N6226,N6227,N6228,N6229,N6230,N6231,N6232,N6235,N6236,N6239,N6240,N6241,N6242,N6243,N6246,N6249,N6252,N6255,N6256,N6257,N6258,N6259,N6260,N6261,N6262,N6263,N6266,N6540,N6541,N6542,N6543,N6544,N6545,N6546,N6547,N6555,N6556,N6557,N6558,N6559,N6560,N6561,N6569,N6594,N6595,N6596,N6597,N6598,N6599,N6600,N6601,N6602,N6603,N6604,N6605,N6606,N6621,N6622,N6623,N6624,N6625,N6626,N6627,N6628,N6629,N6639,N6640,N6641,N6642,N6643,N6644,N6645,N6646,N6647,N6648,N6649,N6650,N6651,N6652,N6653,N6654,N6655,N6656,N6657,N6658,N6659,N6660,N6661,N6668,N6677,N6678,N6679,N6680,N6681,N6682,N6683,N6684,N6685,N6686,N6687,N6688,N6689,N6690,N6702,N6703,N6704,N6705,N6706,N6707,N6708,N6709,N6710,N6711,N6712,N6729,N6730,N6731,N6732,N6733,N6734,N6735,N6736,N6741,N6742,N6743,N6744,N6751,N6752,N6753,N6754,N6755,N6756,N6757,N6758,N6761,N6762,N6766,N6767,N6768,N6769,N6770,N6771,N6772,N6773,N6774,N6775,N6776,N6777,N6778,N6779,N6780,N6781,N6782,N6783,N6784,N6787,N6788,N6789,N6790,N6791,N6792,N6793,N6794,N6795,N6796,N6797,N6800,N6803,N6806,N6809,N6812,N6815,N6818,N6821,N6824,N6827,N6830,N6833,N6836,N6837,N6838,N6839,N6840,N6841,N6842,N6843,N6844,N6845,N6848,N6849,N6850,N6851,N6852,N6853,N6854,N6855,N6856,N6857,N6858,N6859,N6860,N6861,N6862,N6863,N6864,N6865,N6866,N6867,N6870,N6871,N6872,N6873,N6874,N6875,N6876,N6877,N6878,N6879,N6880,N6881,N6884,N6885,N6886,N6887,N6888,N6889,N6890,N6891,N6892,N6893,N6894,N6901,N6912,N6923,N6929,N6936,N6946,N6957,N6967,N6968,N6969,N6970,N6977,N6988,N6998,N7006,N7020,N7036,N7049,N7055,N7056,N7057,N7060,N7061,N7062,N7063,N7064,N7065,N7066,N7067,N7068,N7073,N7077,N7080,N7086,N7091,N7095,N7098,N7099,N7100,N7103,N7104,N7105,N7106,N7107,N7114,N7125,N7136,N7142,N7149,N7159,N7170,N7180,N7187,N7188,N7191,N7194,N7198,N7202,N7205,N7209,N7213,N7216,N7219,N7222,N7229,N7240,N7250,N7258,N7272,N7288,N7301,N7307,N7314,N7318,N7322,N7325,N7328,N7331,N7334,N7337,N7340,N7343,N7346,N7351,N7355,N7358,N7364,N7369,N7373,N7376,N7377,N7378,N7381,N7384,N7387,N7391,N7394,N7398,N7402,N7405,N7408,N7411,N7414,N7417,N7420,N7423,N7426,N7429,N7432,N7435,N7438,N7441,N7444,N7447,N7450,N7453,N7456,N7459,N7462,N7465,N7468,N7471,N7474,N7477,N7478,N7479,N7482,N7485,N7488,N7491,N7494,N7497,N7500,N7503,N7506,N7509,N7512,N7515,N7518,N7521,N7524,N7527,N7530,N7533,N7536,N7539,N7542,N7545,N7548,N7551,N7552,N7553,N7556,N7557,N7558,N7559,N7560,N7563,N7566,N7569,N7572,N7573,N7574,N7577,N7580,N7581,N7582,N7585,N7588,N7591,N7609,N7613,N7620,N7649,N7650,N7655,N7659,N7668,N7671,N7744,N7822,N7825,N7826,N7852,N8114,N8117,N8131,N8134,N8144,N8145,N8146,N8156,N8166,N8169,N8183,N8186,N8196,N8200,N8204,N8208,N8216,N8217,N8218,N8219,N8232,N8233,N8242,N8243,N8244,N8245,N8246,N8247,N8248,N8249,N8250,N8251,N8252,N8253,N8254,N8260,N8261,N8262,N8269,N8274,N8275,N8276,N8277,N8278,N8279,N8280,N8281,N8282,N8283,N8284,N8285,N8288,N8294,N8295,N8296,N8297,N8298,N8307,N8315,N8317,N8319,N8321,N8322,N8323,N8324,N8325,N8326,N8333,N8337,N8338,N8339,N8340,N8341,N8342,N8343,N8344,N8345,N8346,N8347,N8348,N8349,N8350,N8351,N8352,N8353,N8354,N8355,N8356,N8357,N8358,N8365,N8369,N8370,N8371,N8372,N8373,N8374,N8375,N8376,N8377,N8378,N8379,N8380,N8381,N8382,N8383,N8384,N8385,N8386,N8387,N8388,N8389,N8390,N8391,N8392,N8393,N8394,N8404,N8405,N8409,N8410,N8411,N8412,N8415,N8416,N8417,N8418,N8421,N8430,N8433,N8434,N8435,N8436,N8437,N8438,N8439,N8440,N8441,N8442,N8443,N8444,N8447,N8448,N8449,N8450,N8451,N8452,N8453,N8454,N8455,N8456,N8457,N8460,N8463,N8466,N8469,N8470,N8471,N8474,N8477,N8480,N8483,N8484,N8485,N8488,N8489,N8490,N8491,N8492,N8493,N8494,N8495,N8496,N8497,N8500,N8501,N8502,N8503,N8504,N8505,N8506,N8507,N8508,N8509,N8510,N8511,N8512,N8513,N8514,N8515,N8516,N8517,N8518,N8519,N8522,N8525,N8528,N8531,N8534,N8537,N8538,N8539,N8540,N8541,N8545,N8546,N8547,N8548,N8551,N8552,N8553,N8554,N8555,N8558,N8561,N8564,N8565,N8566,N8569,N8572,N8575,N8578,N8579,N8580,N8583,N8586,N8589,N8592,N8595,N8598,N8601,N8604,N8607,N8608,N8609,N8610,N8615,N8616,N8617,N8618,N8619,N8624,N8625,N8626,N8627,N8632,N8633,N8634,N8637,N8638,N8639,N8644,N8645,N8646,N8647,N8648,N8653,N8654,N8655,N8660,N8663,N8666,N8669,N8672,N8675,N8678,N8681,N8684,N8687,N8690,N8693,N8696,N8699,N8702,N8705,N8708,N8711,N8714,N8717,N8718,N8721,N8724,N8727,N8730,N8733,N8734,N8735,N8738,N8741,N8744,N8747,N8750,N8753,N8754,N8755,N8756,N8757,N8760,N8763,N8766,N8769,N8772,N8775,N8778,N8781,N8784,N8787,N8790,N8793,N8796,N8799,N8802,N8805,N8808,N8811,N8814,N8815,N8816,N8817,N8818,N8840,N8857,N8861,N8862,N8863,N8864,N8865,N8866,N8871,N8874,N8878,N8879,N8880,N8881,N8882,N8883,N8884,N8885,N8886,N8887,N8888,N8898,N8902,N8920,N8924,N8927,N8931,N8943,N8950,N8956,N8959,N8960,N8963,N8966,N8991,N8992,N8995,N8996,N9001,N9005,N9024,N9025,N9029,N9035,N9053,N9054,N9064,N9065,N9066,N9067,N9068,N9071,N9072,N9073,N9074,N9077,N9079,N9082,N9083,N9086,N9087,N9088,N9089,N9092,N9093,N9094,N9095,N9098,N9099,N9103,N9107,N9111,N9117,N9127,N9146,N9149,N9159,N9160,N9161,N9165,N9169,N9173,N9179,N9180,N9181,N9182,N9183,N9193,N9203,N9206,N9220,N9223,N9234,N9235,N9236,N9237,N9238,N9242,N9243,N9244,N9245,N9246,N9247,N9248,N9249,N9250,N9251,N9252,N9256,N9257,N9258,N9259,N9260,N9261,N9262,N9265,N9268,N9271,N9272,N9273,N9274,N9275,N9276,N9280,N9285,N9286,N9287,N9288,N9290,N9292,N9294,N9296,N9297,N9298,N9299,N9300,N9301,N9307,N9314,N9315,N9318,N9319,N9320,N9321,N9322,N9323,N9324,N9326,N9332,N9339,N9344,N9352,N9354,N9356,N9358,N9359,N9360,N9361,N9362,N9363,N9364,N9365,N9366,N9367,N9368,N9369,N9370,N9371,N9372,N9375,N9381,N9382,N9383,N9384,N9385,N9392,N9393,N9394,N9395,N9396,N9397,N9398,N9399,N9400,N9401,N9402,N9407,N9408,N9412,N9413,N9414,N9415,N9416,N9417,N9418,N9419,N9420,N9421,N9422,N9423,N9426,N9429,N9432,N9435,N9442,N9445,N9454,N9455,N9456,N9459,N9460,N9461,N9462,N9465,N9466,N9467,N9468,N9473,N9476,N9477,N9478,N9485,N9488,N9493,N9494,N9495,N9498,N9499,N9500,N9505,N9506,N9507,N9508,N9509,N9514,N9515,N9516,N9517,N9520,N9526,N9531,N9539,N9540,N9541,N9543,N9551,N9555,N9556,N9557,N9560,N9561,N9562,N9563,N9564,N9565,N9566,N9567,N9568,N9569,N9570,N9571,N9575,N9579,N9581,N9582,N9585,N9591,N9592,N9593,N9594,N9595,N9596,N9597,N9598,N9599,N9600,N9601,N9602,N9603,N9604,N9605,N9608,N9611,N9612,N9613,N9614,N9615,N9616,N9617,N9618,N9621,N9622,N9623,N9624,N9626,N9629,N9632,N9635,N9642,N9645,N9646,N9649,N9650,N9653,N9656,N9659,N9660,N9661,N9662,N9663,N9666,N9667,N9670,N9671,N9674,N9675,N9678,N9679,N9682,N9685,N9690,N9691,N9692,N9695,N9698,N9702,N9707,N9710,N9711,N9714,N9715,N9716,N9717,N9720,N9721,N9722,N9723,N9726,N9727,N9732,N9733,N9734,N9735,N9736,N9737,N9738,N9739,N9740,N9741,N9742,N9754,N9758,N9762,N9763,N9764,N9765,N9766,N9767,N9768,N9769,N9773,N9774,N9775,N9779,N9784,N9785,N9786,N9790,N9791,N9795,N9796,N9797,N9798,N9799,N9800,N9801,N9802,N9803,N9805,N9806,N9809,N9813,N9814,N9815,N9816,N9817,N9820,N9825,N9826,N9827,N9828,N9829,N9830,N9835,N9836,N9837,N9838,N9846,N9847,N9862,N9863,N9866,N9873,N9876,N9890,N9891,N9892,N9893,N9894,N9895,N9896,N9897,N9898,N9899,N9900,N9901,N9902,N9903,N9904,N9905,N9906,N9907,N9908,N9909,N9910,N9911,N9917,N9923,N9924,N9925,N9932,N9935,N9938,N9939,N9945,N9946,N9947,N9948,N9949,N9953,N9954,N9955,N9956,N9957,N9958,N9959,N9960,N9961,N9964,N9967,N9968,N9969,N9970,N9971,N9972,N9973,N9974,N9975,N9976,N9977,N9978,N9979,N9982,N9983,N9986,N9989,N9992,N9995,N9996,N9997,N9998,N9999,N10002,N10003,N10006,N10007,N10010,N10013,N10014,N10015,N10016,N10017,N10018,N10019,N10020,N10021,N10022,N10023,N10024,N10026,N10028,N10032,N10033,N10034,N10035,N10036,N10037,N10038,N10039,N10040,N10041,N10042,N10043,N10050,N10053,N10054,N10055,N10056,N10057,N10058,N10059,N10060,N10061,N10062,N10067,N10070,N10073,N10076,N10077,N10082,N10083,N10084,N10085,N10086,N10093,N10094,N10105,N10106,N10107,N10108,N10113,N10114,N10115,N10116,N10119,N10124,N10130,N10131,N10132,N10133,N10134,N10135,N10136,N10137,N10138,N10139,N10140,N10141,N10148,N10155,N10156,N10157,N10158,N10159,N10160,N10161,N10162,N10163,N10164,N10165,N10170,N10173,N10176,N10177,N10178,N10179,N10180,N10183,N10186,N10189,N10192,N10195,N10196,N10197,N10200,N10203,N10204,N10205,N10206,N10212,N10213,N10230,N10231,N10232,N10233,N10234,N10237,N10238,N10239,N10240,N10241,N10242,N10247,N10248,N10259,N10264,N10265,N10266,N10267,N10268,N10269,N10270,N10271,N10272,N10273,N10278,N10279,N10280,N10281,N10282,N10283,N10287,N10288,N10289,N10290,N10291,N10292,N10293,N10294,N10295,N10296,N10299,N10300,N10301,N10306,N10307,N10308,N10311,N10314,N10315,N10316,N10317,N10318,N10321,N10324,N10325,N10326,N10327,N10328,N10329,N10330,N10331,N10332,N10333,N10334,N10337,N10338,N10339,N10340,N10341,N10344,N10354,N10357,N10360,N10367,N10375,N10381,N10388,N10391,N10399,N10402,N10406,N10409,N10412,N10415,N10419,N10422,N10425,N10428,N10431,N10432,N10437,N10438,N10439,N10440,N10441,N10444,N10445,N10450,N10451,N10455,N10456,N10465,N10466,N10479,N10497,N10509,N10512,N10515,N10516,N10517,N10518,N10519,N10522,N10525,N10528,N10531,N10534,N10535,N10536,N10539,N10542,N10543,N10544,N10545,N10546,N10547,N10548,N10549,N10550,N10551,N10552,N10553,N10554,N10555,N10556,N10557,N10558,N10559,N10560,N10561,N10562,N10563,N10564,N10565,N10566,N10567,N10568,N10569,N10570,N10571,N10572,N10573,N10577,N10581,N10582,N10583,N10587,N10588,N10589,N10594,N10595,N10596,N10597,N10598,N10602,N10609,N10610,N10621,N10626,N10627,N10629,N10631,N10637,N10638,N10639,N10640,N10642,N10643,N10644,N10645,N10647,N10648,N10649,N10652,N10659,N10662,N10665,N10668,N10671,N10672,N10673,N10674,N10675,N10678,N10681,N10682,N10683,N10684,N10685,N10686,N10687,N10688,N10689,N10690,N10691,N10694,N10695,N10696,N10697,N10698,N10701,N10705,N10707,N10708,N10709,N10710,N10719,N10720,N10730,N10731,N10737,N10738,N10739,N10746,N10747,N10748,N10749,N10750,N10753,N10754,N10764,N10765,N10766,N10767,N10768,N10769,N10770,N10771,N10772,N10773,N10774,N10775,N10776,N10778,N10781,N10784,N10789,N10792,N10796,N10797,N10798,N10799,N10800,N10803,N10806,N10809,N10812,N10815,N10816,N10817,N10820,N10823,N10824,N10825,N10826,N10832,N10833,N10834,N10835,N10836,N10845,N10846,N10857,N10862,N10863,N10864,N10865,N10866,N10867,N10872,N10873,N10874,N10875,N10876,N10879,N10882,N10883,N10884,N10885,N10886,N10887,N10888,N10889,N10890,N10891,N10892,N10895,N10896,N10897,N10898,N10899,N10902,N10909,N10910,N10915,N10916,N10917,N10918,N10919,N10922,N10923,N10928,N10931,N10934,N10935,N10936,N10937,N10938,N10941,N10944,N10947,N10950,N10953,N10954,N10955,N10958,N10961,N10962,N10963,N10964,N10969,N10970,N10981,N10986,N10987,N10988,N10989,N10990,N10991,N10992,N10995,N10998,N10999,N11000,N11001,N11002,N11003,N11004,N11005,N11006,N11007,N11008,N11011,N11012,N11013,N11014,N11015,N11018,N11023,N11024,N11027,N11028,N11029,N11030,N11031,N11034,N11035,N11040,N11041,N11042,N11043,N11044,N11047,N11050,N11053,N11056,N11059,N11062,N11065,N11066,N11067,N11070,N11073,N11074,N11075,N11076,N11077,N11078,N11095,N11098,N11099,N11100,N11103,N11106,N11107,N11108,N11109,N11110,N11111,N11112,N11113,N11114,N11115,N11116,N11117,N11118,N11119,N11120,N11121,N11122,N11123,N11124,N11127,N11130,N11137,N11138,N11139,N11140,N11141,N11142,N11143,N11144,N11145,N11152,N11153,N11154,N11155,N11156,N11159,N11162,N11165,N11168,N11171,N11174,N11177,N11180,N11183,N11184,N11185,N11186,N11187,N11188,N11205,N11210,N11211,N11212,N11213,N11214,N11215,N11216,N11217,N11218,N11219,N11220,N11222,N11223,N11224,N11225,N11226,N11227,N11228,N11229,N11231,N11232,N11233,N11236,N11239,N11242,N11243,N11244,N11245,N11246,N11250,N11252,N11257,N11260,N11261,N11262,N11263,N11264,N11265,N11267,N11268,N11269,N11270,N11272,N11277,N11278,N11279,N11280,N11282,N11283,N11284,N11285,N11286,N11288,N11289,N11290,N11291,N11292,N11293,N11294,N11295,N11296,N11297,N11298,N11299,N11302,N11307,N11308,N11309,N11312,N11313,N11314,N11315,N11316,N11317,N11320,N11321,N11323,N11327,N11328,N11329,N11331,N11335,N11336,N11337,N11338,N11339,N11341;
BUFX1 BUFF1_1 (.Y(N387),.A(N1));
BUFX1 BUFF1_2 (.Y(N388),.A(N1));
INVX1 NOT1_3 (.Y(N467),.A(N57));
AND2X1 AND2_4 (.Y(N469),.A(N134),.B(N133));
BUFX1 BUFF1_5 (.Y(N478),.A(N248));
BUFX1 BUFF1_6 (.Y(N482),.A(N254));
BUFX1 BUFF1_7 (.Y(N484),.A(N257));
BUFX1 BUFF1_8 (.Y(N486),.A(N260));
BUFX1 BUFF1_9 (.Y(N489),.A(N263));
BUFX1 BUFF1_10 (.Y(N492),.A(N267));
AND2X1 AND_tmp1 (.Y(ttmp1),.A(N188),.B(N199));
AND2X1 AND_tmp2 (.Y(ttmp2),.A(N162),.B(ttmp1));
AND2X1 AND_tmp3 (.Y(N494),.A(N172),.B(ttmp2));
BUFX1 BUFF1_12 (.Y(N501),.A(N274));
BUFX1 BUFF1_13 (.Y(N505),.A(N280));
BUFX1 BUFF1_14 (.Y(N507),.A(N283));
BUFX1 BUFF1_15 (.Y(N509),.A(N286));
BUFX1 BUFF1_16 (.Y(N511),.A(N289));
BUFX1 BUFF1_17 (.Y(N513),.A(N293));
BUFX1 BUFF1_18 (.Y(N515),.A(N296));
BUFX1 BUFF1_19 (.Y(N517),.A(N299));
BUFX1 BUFF1_20 (.Y(N519),.A(N303));
AND2X1 AND_tmp4 (.Y(ttmp4),.A(N228),.B(N240));
AND2X1 AND_tmp5 (.Y(ttmp5),.A(N150),.B(ttmp4));
AND2X1 AND_tmp6 (.Y(N528),.A(N184),.B(ttmp5));
BUFX1 BUFF1_22 (.Y(N535),.A(N307));
BUFX1 BUFF1_23 (.Y(N537),.A(N310));
BUFX1 BUFF1_24 (.Y(N539),.A(N313));
BUFX1 BUFF1_25 (.Y(N541),.A(N316));
BUFX1 BUFF1_26 (.Y(N543),.A(N319));
BUFX1 BUFF1_27 (.Y(N545),.A(N322));
BUFX1 BUFF1_28 (.Y(N547),.A(N325));
BUFX1 BUFF1_29 (.Y(N549),.A(N328));
BUFX1 BUFF1_30 (.Y(N551),.A(N331));
BUFX1 BUFF1_31 (.Y(N553),.A(N334));
BUFX1 BUFF1_32 (.Y(N556),.A(N337));
BUFX1 BUFF1_33 (.Y(N559),.A(N343));
BUFX1 BUFF1_34 (.Y(N561),.A(N346));
BUFX1 BUFF1_35 (.Y(N563),.A(N349));
BUFX1 BUFF1_36 (.Y(N565),.A(N352));
BUFX1 BUFF1_37 (.Y(N567),.A(N355));
BUFX1 BUFF1_38 (.Y(N569),.A(N358));
BUFX1 BUFF1_39 (.Y(N571),.A(N361));
BUFX1 BUFF1_40 (.Y(N573),.A(N364));
AND2X1 AND_tmp7 (.Y(ttmp7),.A(N185),.B(N186));
AND2X1 AND_tmp8 (.Y(ttmp8),.A(N183),.B(ttmp7));
AND2X1 AND_tmp9 (.Y(N575),.A(N182),.B(ttmp8));
AND2X1 AND_tmp10 (.Y(ttmp10),.A(N218),.B(N230));
AND2X1 AND_tmp11 (.Y(ttmp11),.A(N210),.B(ttmp10));
AND2X1 AND_tmp12 (.Y(N578),.A(N152),.B(ttmp11));
INVX1 NOT1_43 (.Y(N582),.A(N15));
INVX1 NOT1_44 (.Y(N585),.A(N5));
BUFX1 BUFF1_45 (.Y(N590),.A(N1));
INVX1 NOT1_46 (.Y(N593),.A(N5));
INVX1 NOT1_47 (.Y(N596),.A(N5));
INVX1 NOT1_48 (.Y(N599),.A(N289));
INVX1 NOT1_49 (.Y(N604),.A(N299));
INVX1 NOT1_50 (.Y(N609),.A(N303));
BUFX1 BUFF1_51 (.Y(N614),.A(N38));
BUFX1 BUFF1_52 (.Y(N625),.A(N15));
NAND2X1 NAND2_53 (.Y(N628),.A(N12),.B(N9));
NAND2X1 NAND2_54 (.Y(N632),.A(N12),.B(N9));
BUFX1 BUFF1_55 (.Y(N636),.A(N38));
INVX1 NOT1_56 (.Y(N641),.A(N245));
INVX1 NOT1_57 (.Y(N642),.A(N248));
BUFX1 BUFF1_58 (.Y(N643),.A(N251));
INVX1 NOT1_59 (.Y(N644),.A(N251));
INVX1 NOT1_60 (.Y(N651),.A(N254));
BUFX1 BUFF1_61 (.Y(N657),.A(N106));
INVX1 NOT1_62 (.Y(N660),.A(N257));
INVX1 NOT1_63 (.Y(N666),.A(N260));
INVX1 NOT1_64 (.Y(N672),.A(N263));
INVX1 NOT1_65 (.Y(N673),.A(N267));
INVX1 NOT1_66 (.Y(N674),.A(N106));
BUFX1 BUFF1_67 (.Y(N676),.A(N18));
BUFX1 BUFF1_68 (.Y(N682),.A(N18));
AND2X1 AND2_69 (.Y(N688),.A(N382),.B(N263));
BUFX1 BUFF1_70 (.Y(N689),.A(N18));
INVX1 NOT1_71 (.Y(N695),.A(N18));
NAND2X1 NAND2_72 (.Y(N700),.A(N382),.B(N267));
INVX1 NOT1_73 (.Y(N705),.A(N271));
INVX1 NOT1_74 (.Y(N706),.A(N274));
BUFX1 BUFF1_75 (.Y(N707),.A(N277));
INVX1 NOT1_76 (.Y(N708),.A(N277));
INVX1 NOT1_77 (.Y(N715),.A(N280));
INVX1 NOT1_78 (.Y(N721),.A(N283));
INVX1 NOT1_79 (.Y(N727),.A(N286));
INVX1 NOT1_80 (.Y(N733),.A(N289));
INVX1 NOT1_81 (.Y(N734),.A(N293));
INVX1 NOT1_82 (.Y(N742),.A(N296));
INVX1 NOT1_83 (.Y(N748),.A(N299));
INVX1 NOT1_84 (.Y(N749),.A(N303));
BUFX1 BUFF1_85 (.Y(N750),.A(N367));
INVX1 NOT1_86 (.Y(N758),.A(N307));
INVX1 NOT1_87 (.Y(N759),.A(N310));
INVX1 NOT1_88 (.Y(N762),.A(N313));
INVX1 NOT1_89 (.Y(N768),.A(N316));
INVX1 NOT1_90 (.Y(N774),.A(N319));
INVX1 NOT1_91 (.Y(N780),.A(N322));
INVX1 NOT1_92 (.Y(N786),.A(N325));
INVX1 NOT1_93 (.Y(N794),.A(N328));
INVX1 NOT1_94 (.Y(N800),.A(N331));
INVX1 NOT1_95 (.Y(N806),.A(N334));
INVX1 NOT1_96 (.Y(N812),.A(N337));
BUFX1 BUFF1_97 (.Y(N813),.A(N340));
INVX1 NOT1_98 (.Y(N814),.A(N340));
INVX1 NOT1_99 (.Y(N821),.A(N343));
INVX1 NOT1_100 (.Y(N827),.A(N346));
INVX1 NOT1_101 (.Y(N833),.A(N349));
INVX1 NOT1_102 (.Y(N839),.A(N352));
INVX1 NOT1_103 (.Y(N845),.A(N355));
INVX1 NOT1_104 (.Y(N853),.A(N358));
INVX1 NOT1_105 (.Y(N859),.A(N361));
INVX1 NOT1_106 (.Y(N865),.A(N364));
BUFX1 BUFF1_107 (.Y(N871),.A(N367));
NAND2X1 NAND2_108 (.Y(N881),.A(N467),.B(N585));
INVX1 NOT1_109 (.Y(N882),.A(N528));
INVX1 NOT1_110 (.Y(N883),.A(N578));
INVX1 NOT1_111 (.Y(N884),.A(N575));
INVX1 NOT1_112 (.Y(N885),.A(N494));
AND2X1 AND2_113 (.Y(N886),.A(N528),.B(N578));
AND2X1 AND2_114 (.Y(N887),.A(N575),.B(N494));
BUFX1 BUFF1_115 (.Y(N889),.A(N590));
BUFX1 BUFF1_116 (.Y(N945),.A(N657));
INVX1 NOT1_117 (.Y(N957),.A(N688));
AND2X1 AND2_118 (.Y(N1028),.A(N382),.B(N641));
NAND2X1 NAND2_119 (.Y(N1029),.A(N382),.B(N705));
AND2X1 AND2_120 (.Y(N1109),.A(N469),.B(N596));
NAND2X1 NAND2_121 (.Y(N1110),.A(N242),.B(N593));
INVX1 NOT1_122 (.Y(N1111),.A(N625));
NAND2X1 NAND2_123 (.Y(N1112),.A(N242),.B(N593));
NAND2X1 NAND2_124 (.Y(N1113),.A(N469),.B(N596));
INVX1 NOT1_125 (.Y(N1114),.A(N625));
INVX1 NOT1_126 (.Y(N1115),.A(N871));
BUFX1 BUFF1_127 (.Y(N1116),.A(N590));
BUFX1 BUFF1_128 (.Y(N1119),.A(N628));
BUFX1 BUFF1_129 (.Y(N1125),.A(N682));
BUFX1 BUFF1_130 (.Y(N1132),.A(N628));
BUFX1 BUFF1_131 (.Y(N1136),.A(N682));
BUFX1 BUFF1_132 (.Y(N1141),.A(N628));
BUFX1 BUFF1_133 (.Y(N1147),.A(N682));
BUFX1 BUFF1_134 (.Y(N1154),.A(N632));
BUFX1 BUFF1_135 (.Y(N1160),.A(N676));
AND2X1 AND2_136 (.Y(N1167),.A(N700),.B(N614));
AND2X1 AND2_137 (.Y(N1174),.A(N700),.B(N614));
BUFX1 BUFF1_138 (.Y(N1175),.A(N682));
BUFX1 BUFF1_139 (.Y(N1182),.A(N676));
INVX1 NOT1_140 (.Y(N1189),.A(N657));
INVX1 NOT1_141 (.Y(N1194),.A(N676));
INVX1 NOT1_142 (.Y(N1199),.A(N682));
INVX1 NOT1_143 (.Y(N1206),.A(N689));
BUFX1 BUFF1_144 (.Y(N1211),.A(N695));
INVX1 NOT1_145 (.Y(N1218),.A(N750));
INVX1 NOT1_146 (.Y(N1222),.A(N1028));
BUFX1 BUFF1_147 (.Y(N1227),.A(N632));
BUFX1 BUFF1_148 (.Y(N1233),.A(N676));
BUFX1 BUFF1_149 (.Y(N1240),.A(N632));
BUFX1 BUFF1_150 (.Y(N1244),.A(N676));
BUFX1 BUFF1_151 (.Y(N1249),.A(N689));
BUFX1 BUFF1_152 (.Y(N1256),.A(N689));
BUFX1 BUFF1_153 (.Y(N1263),.A(N695));
BUFX1 BUFF1_154 (.Y(N1270),.A(N689));
BUFX1 BUFF1_155 (.Y(N1277),.A(N689));
BUFX1 BUFF1_156 (.Y(N1284),.A(N700));
BUFX1 BUFF1_157 (.Y(N1287),.A(N614));
BUFX1 BUFF1_158 (.Y(N1290),.A(N666));
BUFX1 BUFF1_159 (.Y(N1293),.A(N660));
BUFX1 BUFF1_160 (.Y(N1296),.A(N651));
BUFX1 BUFF1_161 (.Y(N1299),.A(N614));
BUFX1 BUFF1_162 (.Y(N1302),.A(N644));
BUFX1 BUFF1_163 (.Y(N1305),.A(N700));
BUFX1 BUFF1_164 (.Y(N1308),.A(N614));
BUFX1 BUFF1_165 (.Y(N1311),.A(N614));
BUFX1 BUFF1_166 (.Y(N1314),.A(N666));
BUFX1 BUFF1_167 (.Y(N1317),.A(N660));
BUFX1 BUFF1_168 (.Y(N1320),.A(N651));
BUFX1 BUFF1_169 (.Y(N1323),.A(N644));
BUFX1 BUFF1_170 (.Y(N1326),.A(N609));
BUFX1 BUFF1_171 (.Y(N1329),.A(N604));
BUFX1 BUFF1_172 (.Y(N1332),.A(N742));
BUFX1 BUFF1_173 (.Y(N1335),.A(N599));
BUFX1 BUFF1_174 (.Y(N1338),.A(N727));
BUFX1 BUFF1_175 (.Y(N1341),.A(N721));
BUFX1 BUFF1_176 (.Y(N1344),.A(N715));
BUFX1 BUFF1_177 (.Y(N1347),.A(N734));
BUFX1 BUFF1_178 (.Y(N1350),.A(N708));
BUFX1 BUFF1_179 (.Y(N1353),.A(N609));
BUFX1 BUFF1_180 (.Y(N1356),.A(N604));
BUFX1 BUFF1_181 (.Y(N1359),.A(N742));
BUFX1 BUFF1_182 (.Y(N1362),.A(N734));
BUFX1 BUFF1_183 (.Y(N1365),.A(N599));
BUFX1 BUFF1_184 (.Y(N1368),.A(N727));
BUFX1 BUFF1_185 (.Y(N1371),.A(N721));
BUFX1 BUFF1_186 (.Y(N1374),.A(N715));
BUFX1 BUFF1_187 (.Y(N1377),.A(N708));
BUFX1 BUFF1_188 (.Y(N1380),.A(N806));
BUFX1 BUFF1_189 (.Y(N1383),.A(N800));
BUFX1 BUFF1_190 (.Y(N1386),.A(N794));
BUFX1 BUFF1_191 (.Y(N1389),.A(N786));
BUFX1 BUFF1_192 (.Y(N1392),.A(N780));
BUFX1 BUFF1_193 (.Y(N1395),.A(N774));
BUFX1 BUFF1_194 (.Y(N1398),.A(N768));
BUFX1 BUFF1_195 (.Y(N1401),.A(N762));
BUFX1 BUFF1_196 (.Y(N1404),.A(N806));
BUFX1 BUFF1_197 (.Y(N1407),.A(N800));
BUFX1 BUFF1_198 (.Y(N1410),.A(N794));
BUFX1 BUFF1_199 (.Y(N1413),.A(N780));
BUFX1 BUFF1_200 (.Y(N1416),.A(N774));
BUFX1 BUFF1_201 (.Y(N1419),.A(N768));
BUFX1 BUFF1_202 (.Y(N1422),.A(N762));
BUFX1 BUFF1_203 (.Y(N1425),.A(N786));
BUFX1 BUFF1_204 (.Y(N1428),.A(N636));
BUFX1 BUFF1_205 (.Y(N1431),.A(N636));
BUFX1 BUFF1_206 (.Y(N1434),.A(N865));
BUFX1 BUFF1_207 (.Y(N1437),.A(N859));
BUFX1 BUFF1_208 (.Y(N1440),.A(N853));
BUFX1 BUFF1_209 (.Y(N1443),.A(N845));
BUFX1 BUFF1_210 (.Y(N1446),.A(N839));
BUFX1 BUFF1_211 (.Y(N1449),.A(N833));
BUFX1 BUFF1_212 (.Y(N1452),.A(N827));
BUFX1 BUFF1_213 (.Y(N1455),.A(N821));
BUFX1 BUFF1_214 (.Y(N1458),.A(N814));
BUFX1 BUFF1_215 (.Y(N1461),.A(N865));
BUFX1 BUFF1_216 (.Y(N1464),.A(N859));
BUFX1 BUFF1_217 (.Y(N1467),.A(N853));
BUFX1 BUFF1_218 (.Y(N1470),.A(N839));
BUFX1 BUFF1_219 (.Y(N1473),.A(N833));
BUFX1 BUFF1_220 (.Y(N1476),.A(N827));
BUFX1 BUFF1_221 (.Y(N1479),.A(N821));
BUFX1 BUFF1_222 (.Y(N1482),.A(N845));
BUFX1 BUFF1_223 (.Y(N1485),.A(N814));
INVX1 NOT1_224 (.Y(N1489),.A(N1109));
BUFX1 BUFF1_225 (.Y(N1490),.A(N1116));
AND2X1 AND2_226 (.Y(N1537),.A(N957),.B(N614));
AND2X1 AND2_227 (.Y(N1551),.A(N614),.B(N957));
AND2X1 AND2_228 (.Y(N1649),.A(N1029),.B(N636));
BUFX1 BUFF1_229 (.Y(N1703),.A(N957));
NOR2X1 NOR2_230 (.Y(N1708),.A(N957),.B(N614));
BUFX1 BUFF1_231 (.Y(N1713),.A(N957));
NOR2X1 NOR2_232 (.Y(N1721),.A(N614),.B(N957));
BUFX1 BUFF1_233 (.Y(N1758),.A(N1029));
AND2X1 AND2_234 (.Y(N1781),.A(N163),.B(N1116));
AND2X1 AND2_235 (.Y(N1782),.A(N170),.B(N1125));
INVX1 NOT1_236 (.Y(N1783),.A(N1125));
INVX1 NOT1_237 (.Y(N1789),.A(N1136));
AND2X1 AND2_238 (.Y(N1793),.A(N169),.B(N1125));
AND2X1 AND2_239 (.Y(N1794),.A(N168),.B(N1125));
AND2X1 AND2_240 (.Y(N1795),.A(N167),.B(N1125));
AND2X1 AND2_241 (.Y(N1796),.A(N166),.B(N1136));
AND2X1 AND2_242 (.Y(N1797),.A(N165),.B(N1136));
AND2X1 AND2_243 (.Y(N1798),.A(N164),.B(N1136));
INVX1 NOT1_244 (.Y(N1799),.A(N1147));
INVX1 NOT1_245 (.Y(N1805),.A(N1160));
AND2X1 AND2_246 (.Y(N1811),.A(N177),.B(N1147));
AND2X1 AND2_247 (.Y(N1812),.A(N176),.B(N1147));
AND2X1 AND2_248 (.Y(N1813),.A(N175),.B(N1147));
AND2X1 AND2_249 (.Y(N1814),.A(N174),.B(N1147));
AND2X1 AND2_250 (.Y(N1815),.A(N173),.B(N1147));
AND2X1 AND2_251 (.Y(N1816),.A(N157),.B(N1160));
AND2X1 AND2_252 (.Y(N1817),.A(N156),.B(N1160));
AND2X1 AND2_253 (.Y(N1818),.A(N155),.B(N1160));
AND2X1 AND2_254 (.Y(N1819),.A(N154),.B(N1160));
AND2X1 AND2_255 (.Y(N1820),.A(N153),.B(N1160));
INVX1 NOT1_256 (.Y(N1821),.A(N1284));
INVX1 NOT1_257 (.Y(N1822),.A(N1287));
INVX1 NOT1_258 (.Y(N1828),.A(N1290));
INVX1 NOT1_259 (.Y(N1829),.A(N1293));
INVX1 NOT1_260 (.Y(N1830),.A(N1296));
INVX1 NOT1_261 (.Y(N1832),.A(N1299));
INVX1 NOT1_262 (.Y(N1833),.A(N1302));
INVX1 NOT1_263 (.Y(N1834),.A(N1305));
INVX1 NOT1_264 (.Y(N1835),.A(N1308));
INVX1 NOT1_265 (.Y(N1839),.A(N1311));
INVX1 NOT1_266 (.Y(N1840),.A(N1314));
INVX1 NOT1_267 (.Y(N1841),.A(N1317));
INVX1 NOT1_268 (.Y(N1842),.A(N1320));
INVX1 NOT1_269 (.Y(N1843),.A(N1323));
INVX1 NOT1_270 (.Y(N1845),.A(N1175));
INVX1 NOT1_271 (.Y(N1851),.A(N1182));
AND2X1 AND2_272 (.Y(N1857),.A(N181),.B(N1175));
AND2X1 AND2_273 (.Y(N1858),.A(N171),.B(N1175));
AND2X1 AND2_274 (.Y(N1859),.A(N180),.B(N1175));
AND2X1 AND2_275 (.Y(N1860),.A(N179),.B(N1175));
AND2X1 AND2_276 (.Y(N1861),.A(N178),.B(N1175));
AND2X1 AND2_277 (.Y(N1862),.A(N161),.B(N1182));
AND2X1 AND2_278 (.Y(N1863),.A(N151),.B(N1182));
AND2X1 AND2_279 (.Y(N1864),.A(N160),.B(N1182));
AND2X1 AND2_280 (.Y(N1865),.A(N159),.B(N1182));
AND2X1 AND2_281 (.Y(N1866),.A(N158),.B(N1182));
INVX1 NOT1_282 (.Y(N1867),.A(N1326));
INVX1 NOT1_283 (.Y(N1868),.A(N1329));
INVX1 NOT1_284 (.Y(N1869),.A(N1332));
INVX1 NOT1_285 (.Y(N1870),.A(N1335));
INVX1 NOT1_286 (.Y(N1871),.A(N1338));
INVX1 NOT1_287 (.Y(N1872),.A(N1341));
INVX1 NOT1_288 (.Y(N1873),.A(N1344));
INVX1 NOT1_289 (.Y(N1874),.A(N1347));
INVX1 NOT1_290 (.Y(N1875),.A(N1350));
INVX1 NOT1_291 (.Y(N1876),.A(N1353));
INVX1 NOT1_292 (.Y(N1877),.A(N1356));
INVX1 NOT1_293 (.Y(N1878),.A(N1359));
INVX1 NOT1_294 (.Y(N1879),.A(N1362));
INVX1 NOT1_295 (.Y(N1880),.A(N1365));
INVX1 NOT1_296 (.Y(N1881),.A(N1368));
INVX1 NOT1_297 (.Y(N1882),.A(N1371));
INVX1 NOT1_298 (.Y(N1883),.A(N1374));
INVX1 NOT1_299 (.Y(N1884),.A(N1377));
BUFX1 BUFF1_300 (.Y(N1885),.A(N1199));
BUFX1 BUFF1_301 (.Y(N1892),.A(N1194));
BUFX1 BUFF1_302 (.Y(N1899),.A(N1199));
BUFX1 BUFF1_303 (.Y(N1906),.A(N1194));
INVX1 NOT1_304 (.Y(N1913),.A(N1211));
BUFX1 BUFF1_305 (.Y(N1919),.A(N1194));
AND2X1 AND2_306 (.Y(N1926),.A(N44),.B(N1211));
AND2X1 AND2_307 (.Y(N1927),.A(N41),.B(N1211));
AND2X1 AND2_308 (.Y(N1928),.A(N29),.B(N1211));
AND2X1 AND2_309 (.Y(N1929),.A(N26),.B(N1211));
AND2X1 AND2_310 (.Y(N1930),.A(N23),.B(N1211));
INVX1 NOT1_311 (.Y(N1931),.A(N1380));
INVX1 NOT1_312 (.Y(N1932),.A(N1383));
INVX1 NOT1_313 (.Y(N1933),.A(N1386));
INVX1 NOT1_314 (.Y(N1934),.A(N1389));
INVX1 NOT1_315 (.Y(N1935),.A(N1392));
INVX1 NOT1_316 (.Y(N1936),.A(N1395));
INVX1 NOT1_317 (.Y(N1937),.A(N1398));
INVX1 NOT1_318 (.Y(N1938),.A(N1401));
INVX1 NOT1_319 (.Y(N1939),.A(N1404));
INVX1 NOT1_320 (.Y(N1940),.A(N1407));
INVX1 NOT1_321 (.Y(N1941),.A(N1410));
INVX1 NOT1_322 (.Y(N1942),.A(N1413));
INVX1 NOT1_323 (.Y(N1943),.A(N1416));
INVX1 NOT1_324 (.Y(N1944),.A(N1419));
INVX1 NOT1_325 (.Y(N1945),.A(N1422));
INVX1 NOT1_326 (.Y(N1946),.A(N1425));
INVX1 NOT1_327 (.Y(N1947),.A(N1233));
INVX1 NOT1_328 (.Y(N1953),.A(N1244));
AND2X1 AND2_329 (.Y(N1957),.A(N209),.B(N1233));
AND2X1 AND2_330 (.Y(N1958),.A(N216),.B(N1233));
AND2X1 AND2_331 (.Y(N1959),.A(N215),.B(N1233));
AND2X1 AND2_332 (.Y(N1960),.A(N214),.B(N1233));
AND2X1 AND2_333 (.Y(N1961),.A(N213),.B(N1244));
AND2X1 AND2_334 (.Y(N1962),.A(N212),.B(N1244));
AND2X1 AND2_335 (.Y(N1963),.A(N211),.B(N1244));
INVX1 NOT1_336 (.Y(N1965),.A(N1428));
AND2X1 AND2_337 (.Y(N1966),.A(N1222),.B(N636));
INVX1 NOT1_338 (.Y(N1967),.A(N1431));
INVX1 NOT1_339 (.Y(N1968),.A(N1434));
INVX1 NOT1_340 (.Y(N1969),.A(N1437));
INVX1 NOT1_341 (.Y(N1970),.A(N1440));
INVX1 NOT1_342 (.Y(N1971),.A(N1443));
INVX1 NOT1_343 (.Y(N1972),.A(N1446));
INVX1 NOT1_344 (.Y(N1973),.A(N1449));
INVX1 NOT1_345 (.Y(N1974),.A(N1452));
INVX1 NOT1_346 (.Y(N1975),.A(N1455));
INVX1 NOT1_347 (.Y(N1976),.A(N1458));
INVX1 NOT1_348 (.Y(N1977),.A(N1249));
INVX1 NOT1_349 (.Y(N1983),.A(N1256));
AND2X1 AND2_350 (.Y(N1989),.A(N642),.B(N1249));
AND2X1 AND2_351 (.Y(N1990),.A(N644),.B(N1249));
AND2X1 AND2_352 (.Y(N1991),.A(N651),.B(N1249));
AND2X1 AND2_353 (.Y(N1992),.A(N674),.B(N1249));
AND2X1 AND2_354 (.Y(N1993),.A(N660),.B(N1249));
AND2X1 AND2_355 (.Y(N1994),.A(N666),.B(N1256));
AND2X1 AND2_356 (.Y(N1995),.A(N672),.B(N1256));
AND2X1 AND2_357 (.Y(N1996),.A(N673),.B(N1256));
INVX1 NOT1_358 (.Y(N1997),.A(N1263));
BUFX1 BUFF1_359 (.Y(N2003),.A(N1194));
AND2X1 AND2_360 (.Y(N2010),.A(N47),.B(N1263));
AND2X1 AND2_361 (.Y(N2011),.A(N35),.B(N1263));
AND2X1 AND2_362 (.Y(N2012),.A(N32),.B(N1263));
AND2X1 AND2_363 (.Y(N2013),.A(N50),.B(N1263));
AND2X1 AND2_364 (.Y(N2014),.A(N66),.B(N1263));
INVX1 NOT1_365 (.Y(N2015),.A(N1461));
INVX1 NOT1_366 (.Y(N2016),.A(N1464));
INVX1 NOT1_367 (.Y(N2017),.A(N1467));
INVX1 NOT1_368 (.Y(N2018),.A(N1470));
INVX1 NOT1_369 (.Y(N2019),.A(N1473));
INVX1 NOT1_370 (.Y(N2020),.A(N1476));
INVX1 NOT1_371 (.Y(N2021),.A(N1479));
INVX1 NOT1_372 (.Y(N2022),.A(N1482));
INVX1 NOT1_373 (.Y(N2023),.A(N1485));
BUFX1 BUFF1_374 (.Y(N2024),.A(N1206));
BUFX1 BUFF1_375 (.Y(N2031),.A(N1206));
BUFX1 BUFF1_376 (.Y(N2038),.A(N1206));
BUFX1 BUFF1_377 (.Y(N2045),.A(N1206));
INVX1 NOT1_378 (.Y(N2052),.A(N1270));
INVX1 NOT1_379 (.Y(N2058),.A(N1277));
AND2X1 AND2_380 (.Y(N2064),.A(N706),.B(N1270));
AND2X1 AND2_381 (.Y(N2065),.A(N708),.B(N1270));
AND2X1 AND2_382 (.Y(N2066),.A(N715),.B(N1270));
AND2X1 AND2_383 (.Y(N2067),.A(N721),.B(N1270));
AND2X1 AND2_384 (.Y(N2068),.A(N727),.B(N1270));
AND2X1 AND2_385 (.Y(N2069),.A(N733),.B(N1277));
AND2X1 AND2_386 (.Y(N2070),.A(N734),.B(N1277));
AND2X1 AND2_387 (.Y(N2071),.A(N742),.B(N1277));
AND2X1 AND2_388 (.Y(N2072),.A(N748),.B(N1277));
AND2X1 AND2_389 (.Y(N2073),.A(N749),.B(N1277));
BUFX1 BUFF1_390 (.Y(N2074),.A(N1189));
BUFX1 BUFF1_391 (.Y(N2081),.A(N1189));
BUFX1 BUFF1_392 (.Y(N2086),.A(N1222));
NAND2X1 NAND2_393 (.Y(N2107),.A(N1287),.B(N1821));
NAND2X1 NAND2_394 (.Y(N2108),.A(N1284),.B(N1822));
INVX1 NOT1_395 (.Y(N2110),.A(N1703));
NAND2X1 NAND2_396 (.Y(N2111),.A(N1703),.B(N1832));
NAND2X1 NAND2_397 (.Y(N2112),.A(N1308),.B(N1834));
NAND2X1 NAND2_398 (.Y(N2113),.A(N1305),.B(N1835));
INVX1 NOT1_399 (.Y(N2114),.A(N1713));
NAND2X1 NAND2_400 (.Y(N2115),.A(N1713),.B(N1839));
INVX1 NOT1_401 (.Y(N2117),.A(N1721));
INVX1 NOT1_402 (.Y(N2171),.A(N1758));
NAND2X1 NAND2_403 (.Y(N2172),.A(N1758),.B(N1965));
INVX1 NOT1_404 (.Y(N2230),.A(N1708));
BUFX1 BUFF1_405 (.Y(N2231),.A(N1537));
BUFX1 BUFF1_406 (.Y(N2235),.A(N1551));
OR2X1 OR2_407 (.Y(N2239),.A(N1783),.B(N1782));
OR2X1 OR2_408 (.Y(N2240),.A(N1783),.B(N1125));
OR2X1 OR2_409 (.Y(N2241),.A(N1783),.B(N1793));
OR2X1 OR2_410 (.Y(N2242),.A(N1783),.B(N1794));
OR2X1 OR2_411 (.Y(N2243),.A(N1783),.B(N1795));
OR2X1 OR2_412 (.Y(N2244),.A(N1789),.B(N1796));
OR2X1 OR2_413 (.Y(N2245),.A(N1789),.B(N1797));
OR2X1 OR2_414 (.Y(N2246),.A(N1789),.B(N1798));
OR2X1 OR2_415 (.Y(N2247),.A(N1799),.B(N1811));
OR2X1 OR2_416 (.Y(N2248),.A(N1799),.B(N1812));
OR2X1 OR2_417 (.Y(N2249),.A(N1799),.B(N1813));
OR2X1 OR2_418 (.Y(N2250),.A(N1799),.B(N1814));
OR2X1 OR2_419 (.Y(N2251),.A(N1799),.B(N1815));
OR2X1 OR2_420 (.Y(N2252),.A(N1805),.B(N1816));
OR2X1 OR2_421 (.Y(N2253),.A(N1805),.B(N1817));
OR2X1 OR2_422 (.Y(N2254),.A(N1805),.B(N1818));
OR2X1 OR2_423 (.Y(N2255),.A(N1805),.B(N1819));
OR2X1 OR2_424 (.Y(N2256),.A(N1805),.B(N1820));
NAND2X1 NAND2_425 (.Y(N2257),.A(N2107),.B(N2108));
INVX1 NOT1_426 (.Y(N2267),.A(N2074));
NAND2X1 NAND2_427 (.Y(N2268),.A(N1299),.B(N2110));
NAND2X1 NAND2_428 (.Y(N2269),.A(N2112),.B(N2113));
NAND2X1 NAND2_429 (.Y(N2274),.A(N1311),.B(N2114));
INVX1 NOT1_430 (.Y(N2275),.A(N2081));
AND2X1 AND2_431 (.Y(N2277),.A(N141),.B(N1845));
AND2X1 AND2_432 (.Y(N2278),.A(N147),.B(N1845));
AND2X1 AND2_433 (.Y(N2279),.A(N138),.B(N1845));
AND2X1 AND2_434 (.Y(N2280),.A(N144),.B(N1845));
AND2X1 AND2_435 (.Y(N2281),.A(N135),.B(N1845));
AND2X1 AND2_436 (.Y(N2282),.A(N141),.B(N1851));
AND2X1 AND2_437 (.Y(N2283),.A(N147),.B(N1851));
AND2X1 AND2_438 (.Y(N2284),.A(N138),.B(N1851));
AND2X1 AND2_439 (.Y(N2285),.A(N144),.B(N1851));
AND2X1 AND2_440 (.Y(N2286),.A(N135),.B(N1851));
INVX1 NOT1_441 (.Y(N2287),.A(N1885));
INVX1 NOT1_442 (.Y(N2293),.A(N1892));
AND2X1 AND2_443 (.Y(N2299),.A(N103),.B(N1885));
AND2X1 AND2_444 (.Y(N2300),.A(N130),.B(N1885));
AND2X1 AND2_445 (.Y(N2301),.A(N127),.B(N1885));
AND2X1 AND2_446 (.Y(N2302),.A(N124),.B(N1885));
AND2X1 AND2_447 (.Y(N2303),.A(N100),.B(N1885));
AND2X1 AND2_448 (.Y(N2304),.A(N103),.B(N1892));
AND2X1 AND2_449 (.Y(N2305),.A(N130),.B(N1892));
AND2X1 AND2_450 (.Y(N2306),.A(N127),.B(N1892));
AND2X1 AND2_451 (.Y(N2307),.A(N124),.B(N1892));
AND2X1 AND2_452 (.Y(N2308),.A(N100),.B(N1892));
INVX1 NOT1_453 (.Y(N2309),.A(N1899));
INVX1 NOT1_454 (.Y(N2315),.A(N1906));
AND2X1 AND2_455 (.Y(N2321),.A(N115),.B(N1899));
AND2X1 AND2_456 (.Y(N2322),.A(N118),.B(N1899));
AND2X1 AND2_457 (.Y(N2323),.A(N97),.B(N1899));
AND2X1 AND2_458 (.Y(N2324),.A(N94),.B(N1899));
AND2X1 AND2_459 (.Y(N2325),.A(N121),.B(N1899));
AND2X1 AND2_460 (.Y(N2326),.A(N115),.B(N1906));
AND2X1 AND2_461 (.Y(N2327),.A(N118),.B(N1906));
AND2X1 AND2_462 (.Y(N2328),.A(N97),.B(N1906));
AND2X1 AND2_463 (.Y(N2329),.A(N94),.B(N1906));
AND2X1 AND2_464 (.Y(N2330),.A(N121),.B(N1906));
INVX1 NOT1_465 (.Y(N2331),.A(N1919));
AND2X1 AND2_466 (.Y(N2337),.A(N208),.B(N1913));
AND2X1 AND2_467 (.Y(N2338),.A(N198),.B(N1913));
AND2X1 AND2_468 (.Y(N2339),.A(N207),.B(N1913));
AND2X1 AND2_469 (.Y(N2340),.A(N206),.B(N1913));
AND2X1 AND2_470 (.Y(N2341),.A(N205),.B(N1913));
AND2X1 AND2_471 (.Y(N2342),.A(N44),.B(N1919));
AND2X1 AND2_472 (.Y(N2343),.A(N41),.B(N1919));
AND2X1 AND2_473 (.Y(N2344),.A(N29),.B(N1919));
AND2X1 AND2_474 (.Y(N2345),.A(N26),.B(N1919));
AND2X1 AND2_475 (.Y(N2346),.A(N23),.B(N1919));
OR2X1 OR2_476 (.Y(N2347),.A(N1947),.B(N1233));
OR2X1 OR2_477 (.Y(N2348),.A(N1947),.B(N1957));
OR2X1 OR2_478 (.Y(N2349),.A(N1947),.B(N1958));
OR2X1 OR2_479 (.Y(N2350),.A(N1947),.B(N1959));
OR2X1 OR2_480 (.Y(N2351),.A(N1947),.B(N1960));
OR2X1 OR2_481 (.Y(N2352),.A(N1953),.B(N1961));
OR2X1 OR2_482 (.Y(N2353),.A(N1953),.B(N1962));
OR2X1 OR2_483 (.Y(N2354),.A(N1953),.B(N1963));
NAND2X1 NAND2_484 (.Y(N2355),.A(N1428),.B(N2171));
INVX1 NOT1_485 (.Y(N2356),.A(N2086));
NAND2X1 NAND2_486 (.Y(N2357),.A(N2086),.B(N1967));
AND2X1 AND2_487 (.Y(N2358),.A(N114),.B(N1977));
AND2X1 AND2_488 (.Y(N2359),.A(N113),.B(N1977));
AND2X1 AND2_489 (.Y(N2360),.A(N111),.B(N1977));
AND2X1 AND2_490 (.Y(N2361),.A(N87),.B(N1977));
AND2X1 AND2_491 (.Y(N2362),.A(N112),.B(N1977));
AND2X1 AND2_492 (.Y(N2363),.A(N88),.B(N1983));
AND2X1 AND2_493 (.Y(N2364),.A(N245),.B(N1983));
AND2X1 AND2_494 (.Y(N2365),.A(N271),.B(N1983));
AND2X1 AND2_495 (.Y(N2366),.A(N759),.B(N1983));
AND2X1 AND2_496 (.Y(N2367),.A(N70),.B(N1983));
INVX1 NOT1_497 (.Y(N2368),.A(N2003));
AND2X1 AND2_498 (.Y(N2374),.A(N193),.B(N1997));
AND2X1 AND2_499 (.Y(N2375),.A(N192),.B(N1997));
AND2X1 AND2_500 (.Y(N2376),.A(N191),.B(N1997));
AND2X1 AND2_501 (.Y(N2377),.A(N190),.B(N1997));
AND2X1 AND2_502 (.Y(N2378),.A(N189),.B(N1997));
AND2X1 AND2_503 (.Y(N2379),.A(N47),.B(N2003));
AND2X1 AND2_504 (.Y(N2380),.A(N35),.B(N2003));
AND2X1 AND2_505 (.Y(N2381),.A(N32),.B(N2003));
AND2X1 AND2_506 (.Y(N2382),.A(N50),.B(N2003));
AND2X1 AND2_507 (.Y(N2383),.A(N66),.B(N2003));
INVX1 NOT1_508 (.Y(N2384),.A(N2024));
INVX1 NOT1_509 (.Y(N2390),.A(N2031));
AND2X1 AND2_510 (.Y(N2396),.A(N58),.B(N2024));
AND2X1 AND2_511 (.Y(N2397),.A(N77),.B(N2024));
AND2X1 AND2_512 (.Y(N2398),.A(N78),.B(N2024));
AND2X1 AND2_513 (.Y(N2399),.A(N59),.B(N2024));
AND2X1 AND2_514 (.Y(N2400),.A(N81),.B(N2024));
AND2X1 AND2_515 (.Y(N2401),.A(N80),.B(N2031));
AND2X1 AND2_516 (.Y(N2402),.A(N79),.B(N2031));
AND2X1 AND2_517 (.Y(N2403),.A(N60),.B(N2031));
AND2X1 AND2_518 (.Y(N2404),.A(N61),.B(N2031));
AND2X1 AND2_519 (.Y(N2405),.A(N62),.B(N2031));
INVX1 NOT1_520 (.Y(N2406),.A(N2038));
INVX1 NOT1_521 (.Y(N2412),.A(N2045));
AND2X1 AND2_522 (.Y(N2418),.A(N69),.B(N2038));
AND2X1 AND2_523 (.Y(N2419),.A(N70),.B(N2038));
AND2X1 AND2_524 (.Y(N2420),.A(N74),.B(N2038));
AND2X1 AND2_525 (.Y(N2421),.A(N76),.B(N2038));
AND2X1 AND2_526 (.Y(N2422),.A(N75),.B(N2038));
AND2X1 AND2_527 (.Y(N2423),.A(N73),.B(N2045));
AND2X1 AND2_528 (.Y(N2424),.A(N53),.B(N2045));
AND2X1 AND2_529 (.Y(N2425),.A(N54),.B(N2045));
AND2X1 AND2_530 (.Y(N2426),.A(N55),.B(N2045));
AND2X1 AND2_531 (.Y(N2427),.A(N56),.B(N2045));
AND2X1 AND2_532 (.Y(N2428),.A(N82),.B(N2052));
AND2X1 AND2_533 (.Y(N2429),.A(N65),.B(N2052));
AND2X1 AND2_534 (.Y(N2430),.A(N83),.B(N2052));
AND2X1 AND2_535 (.Y(N2431),.A(N84),.B(N2052));
AND2X1 AND2_536 (.Y(N2432),.A(N85),.B(N2052));
AND2X1 AND2_537 (.Y(N2433),.A(N64),.B(N2058));
AND2X1 AND2_538 (.Y(N2434),.A(N63),.B(N2058));
AND2X1 AND2_539 (.Y(N2435),.A(N86),.B(N2058));
AND2X1 AND2_540 (.Y(N2436),.A(N109),.B(N2058));
AND2X1 AND2_541 (.Y(N2437),.A(N110),.B(N2058));
AND2X1 AND2_542 (.Y(N2441),.A(N2239),.B(N1119));
AND2X1 AND2_543 (.Y(N2442),.A(N2240),.B(N1119));
AND2X1 AND2_544 (.Y(N2446),.A(N2241),.B(N1119));
AND2X1 AND2_545 (.Y(N2450),.A(N2242),.B(N1119));
AND2X1 AND2_546 (.Y(N2454),.A(N2243),.B(N1119));
AND2X1 AND2_547 (.Y(N2458),.A(N2244),.B(N1132));
AND2X1 AND2_548 (.Y(N2462),.A(N2247),.B(N1141));
AND2X1 AND2_549 (.Y(N2466),.A(N2248),.B(N1141));
AND2X1 AND2_550 (.Y(N2470),.A(N2249),.B(N1141));
AND2X1 AND2_551 (.Y(N2474),.A(N2250),.B(N1141));
AND2X1 AND2_552 (.Y(N2478),.A(N2251),.B(N1141));
AND2X1 AND2_553 (.Y(N2482),.A(N2252),.B(N1154));
AND2X1 AND2_554 (.Y(N2488),.A(N2253),.B(N1154));
AND2X1 AND2_555 (.Y(N2496),.A(N2254),.B(N1154));
AND2X1 AND2_556 (.Y(N2502),.A(N2255),.B(N1154));
AND2X1 AND2_557 (.Y(N2508),.A(N2256),.B(N1154));
NAND2X1 NAND2_558 (.Y(N2523),.A(N2268),.B(N2111));
NAND2X1 NAND2_559 (.Y(N2533),.A(N2274),.B(N2115));
INVX1 NOT1_560 (.Y(N2537),.A(N2235));
OR2X1 OR2_561 (.Y(N2538),.A(N2278),.B(N1858));
OR2X1 OR2_562 (.Y(N2542),.A(N2279),.B(N1859));
OR2X1 OR2_563 (.Y(N2546),.A(N2280),.B(N1860));
OR2X1 OR2_564 (.Y(N2550),.A(N2281),.B(N1861));
OR2X1 OR2_565 (.Y(N2554),.A(N2283),.B(N1863));
OR2X1 OR2_566 (.Y(N2561),.A(N2284),.B(N1864));
OR2X1 OR2_567 (.Y(N2567),.A(N2285),.B(N1865));
OR2X1 OR2_568 (.Y(N2573),.A(N2286),.B(N1866));
OR2X1 OR2_569 (.Y(N2604),.A(N2338),.B(N1927));
OR2X1 OR2_570 (.Y(N2607),.A(N2339),.B(N1928));
OR2X1 OR2_571 (.Y(N2611),.A(N2340),.B(N1929));
OR2X1 OR2_572 (.Y(N2615),.A(N2341),.B(N1930));
AND2X1 AND2_573 (.Y(N2619),.A(N2348),.B(N1227));
AND2X1 AND2_574 (.Y(N2626),.A(N2349),.B(N1227));
AND2X1 AND2_575 (.Y(N2632),.A(N2350),.B(N1227));
AND2X1 AND2_576 (.Y(N2638),.A(N2351),.B(N1227));
AND2X1 AND2_577 (.Y(N2644),.A(N2352),.B(N1240));
NAND2X1 NAND2_578 (.Y(N2650),.A(N2355),.B(N2172));
NAND2X1 NAND2_579 (.Y(N2653),.A(N1431),.B(N2356));
OR2X1 OR2_580 (.Y(N2654),.A(N2359),.B(N1990));
OR2X1 OR2_581 (.Y(N2658),.A(N2360),.B(N1991));
OR2X1 OR2_582 (.Y(N2662),.A(N2361),.B(N1992));
OR2X1 OR2_583 (.Y(N2666),.A(N2362),.B(N1993));
OR2X1 OR2_584 (.Y(N2670),.A(N2363),.B(N1994));
OR2X1 OR2_585 (.Y(N2674),.A(N2366),.B(N1256));
OR2X1 OR2_586 (.Y(N2680),.A(N2367),.B(N1256));
OR2X1 OR2_587 (.Y(N2688),.A(N2374),.B(N2010));
OR2X1 OR2_588 (.Y(N2692),.A(N2375),.B(N2011));
OR2X1 OR2_589 (.Y(N2696),.A(N2376),.B(N2012));
OR2X1 OR2_590 (.Y(N2700),.A(N2377),.B(N2013));
OR2X1 OR2_591 (.Y(N2704),.A(N2378),.B(N2014));
AND2X1 AND2_592 (.Y(N2728),.A(N2347),.B(N1227));
OR2X1 OR2_593 (.Y(N2729),.A(N2429),.B(N2065));
OR2X1 OR2_594 (.Y(N2733),.A(N2430),.B(N2066));
OR2X1 OR2_595 (.Y(N2737),.A(N2431),.B(N2067));
OR2X1 OR2_596 (.Y(N2741),.A(N2432),.B(N2068));
OR2X1 OR2_597 (.Y(N2745),.A(N2433),.B(N2069));
OR2X1 OR2_598 (.Y(N2749),.A(N2434),.B(N2070));
OR2X1 OR2_599 (.Y(N2753),.A(N2435),.B(N2071));
OR2X1 OR2_600 (.Y(N2757),.A(N2436),.B(N2072));
OR2X1 OR2_601 (.Y(N2761),.A(N2437),.B(N2073));
INVX1 NOT1_602 (.Y(N2765),.A(N2231));
AND2X1 AND2_603 (.Y(N2766),.A(N2354),.B(N1240));
AND2X1 AND2_604 (.Y(N2769),.A(N2353),.B(N1240));
AND2X1 AND2_605 (.Y(N2772),.A(N2246),.B(N1132));
AND2X1 AND2_606 (.Y(N2775),.A(N2245),.B(N1132));
OR2X1 OR2_607 (.Y(N2778),.A(N2282),.B(N1862));
OR2X1 OR2_608 (.Y(N2781),.A(N2358),.B(N1989));
OR2X1 OR2_609 (.Y(N2784),.A(N2365),.B(N1996));
OR2X1 OR2_610 (.Y(N2787),.A(N2364),.B(N1995));
OR2X1 OR2_611 (.Y(N2790),.A(N2337),.B(N1926));
OR2X1 OR2_612 (.Y(N2793),.A(N2277),.B(N1857));
OR2X1 OR2_613 (.Y(N2796),.A(N2428),.B(N2064));
AND2X1 AND2_614 (.Y(N2866),.A(N2257),.B(N1537));
AND2X1 AND2_615 (.Y(N2867),.A(N2257),.B(N1537));
AND2X1 AND2_616 (.Y(N2868),.A(N2257),.B(N1537));
AND2X1 AND2_617 (.Y(N2869),.A(N2257),.B(N1537));
AND2X1 AND2_618 (.Y(N2878),.A(N2269),.B(N1551));
AND2X1 AND2_619 (.Y(N2913),.A(N204),.B(N2287));
AND2X1 AND2_620 (.Y(N2914),.A(N203),.B(N2287));
AND2X1 AND2_621 (.Y(N2915),.A(N202),.B(N2287));
AND2X1 AND2_622 (.Y(N2916),.A(N201),.B(N2287));
AND2X1 AND2_623 (.Y(N2917),.A(N200),.B(N2287));
AND2X1 AND2_624 (.Y(N2918),.A(N235),.B(N2293));
AND2X1 AND2_625 (.Y(N2919),.A(N234),.B(N2293));
AND2X1 AND2_626 (.Y(N2920),.A(N233),.B(N2293));
AND2X1 AND2_627 (.Y(N2921),.A(N232),.B(N2293));
AND2X1 AND2_628 (.Y(N2922),.A(N231),.B(N2293));
AND2X1 AND2_629 (.Y(N2923),.A(N197),.B(N2309));
AND2X1 AND2_630 (.Y(N2924),.A(N187),.B(N2309));
AND2X1 AND2_631 (.Y(N2925),.A(N196),.B(N2309));
AND2X1 AND2_632 (.Y(N2926),.A(N195),.B(N2309));
AND2X1 AND2_633 (.Y(N2927),.A(N194),.B(N2309));
AND2X1 AND2_634 (.Y(N2928),.A(N227),.B(N2315));
AND2X1 AND2_635 (.Y(N2929),.A(N217),.B(N2315));
AND2X1 AND2_636 (.Y(N2930),.A(N226),.B(N2315));
AND2X1 AND2_637 (.Y(N2931),.A(N225),.B(N2315));
AND2X1 AND2_638 (.Y(N2932),.A(N224),.B(N2315));
AND2X1 AND2_639 (.Y(N2933),.A(N239),.B(N2331));
AND2X1 AND2_640 (.Y(N2934),.A(N229),.B(N2331));
AND2X1 AND2_641 (.Y(N2935),.A(N238),.B(N2331));
AND2X1 AND2_642 (.Y(N2936),.A(N237),.B(N2331));
AND2X1 AND2_643 (.Y(N2937),.A(N236),.B(N2331));
NAND2X1 NAND2_644 (.Y(N2988),.A(N2653),.B(N2357));
AND2X1 AND2_645 (.Y(N3005),.A(N223),.B(N2368));
AND2X1 AND2_646 (.Y(N3006),.A(N222),.B(N2368));
AND2X1 AND2_647 (.Y(N3007),.A(N221),.B(N2368));
AND2X1 AND2_648 (.Y(N3008),.A(N220),.B(N2368));
AND2X1 AND2_649 (.Y(N3009),.A(N219),.B(N2368));
AND2X1 AND2_650 (.Y(N3020),.A(N812),.B(N2384));
AND2X1 AND2_651 (.Y(N3021),.A(N814),.B(N2384));
AND2X1 AND2_652 (.Y(N3022),.A(N821),.B(N2384));
AND2X1 AND2_653 (.Y(N3023),.A(N827),.B(N2384));
AND2X1 AND2_654 (.Y(N3024),.A(N833),.B(N2384));
AND2X1 AND2_655 (.Y(N3025),.A(N839),.B(N2390));
AND2X1 AND2_656 (.Y(N3026),.A(N845),.B(N2390));
AND2X1 AND2_657 (.Y(N3027),.A(N853),.B(N2390));
AND2X1 AND2_658 (.Y(N3028),.A(N859),.B(N2390));
AND2X1 AND2_659 (.Y(N3029),.A(N865),.B(N2390));
AND2X1 AND2_660 (.Y(N3032),.A(N758),.B(N2406));
AND2X1 AND2_661 (.Y(N3033),.A(N759),.B(N2406));
AND2X1 AND2_662 (.Y(N3034),.A(N762),.B(N2406));
AND2X1 AND2_663 (.Y(N3035),.A(N768),.B(N2406));
AND2X1 AND2_664 (.Y(N3036),.A(N774),.B(N2406));
AND2X1 AND2_665 (.Y(N3037),.A(N780),.B(N2412));
AND2X1 AND2_666 (.Y(N3038),.A(N786),.B(N2412));
AND2X1 AND2_667 (.Y(N3039),.A(N794),.B(N2412));
AND2X1 AND2_668 (.Y(N3040),.A(N800),.B(N2412));
AND2X1 AND2_669 (.Y(N3041),.A(N806),.B(N2412));
BUFX1 BUFF1_670 (.Y(N3061),.A(N2257));
BUFX1 BUFF1_671 (.Y(N3064),.A(N2257));
BUFX1 BUFF1_672 (.Y(N3067),.A(N2269));
BUFX1 BUFF1_673 (.Y(N3070),.A(N2269));
INVX1 NOT1_674 (.Y(N3073),.A(N2728));
INVX1 NOT1_675 (.Y(N3080),.A(N2441));
AND2X1 AND2_676 (.Y(N3096),.A(N666),.B(N2644));
AND2X1 AND2_677 (.Y(N3097),.A(N660),.B(N2638));
AND2X1 AND2_678 (.Y(N3101),.A(N1189),.B(N2632));
AND2X1 AND2_679 (.Y(N3107),.A(N651),.B(N2626));
AND2X1 AND2_680 (.Y(N3114),.A(N644),.B(N2619));
AND2X1 AND2_681 (.Y(N3122),.A(N2523),.B(N2257));
OR2X1 OR2_682 (.Y(N3126),.A(N1167),.B(N2866));
AND2X1 AND2_683 (.Y(N3130),.A(N2523),.B(N2257));
OR2X1 OR2_684 (.Y(N3131),.A(N1167),.B(N2869));
AND2X1 AND2_685 (.Y(N3134),.A(N2523),.B(N2257));
INVX1 NOT1_686 (.Y(N3135),.A(N2533));
AND2X1 AND2_687 (.Y(N3136),.A(N666),.B(N2644));
AND2X1 AND2_688 (.Y(N3137),.A(N660),.B(N2638));
AND2X1 AND2_689 (.Y(N3140),.A(N1189),.B(N2632));
AND2X1 AND2_690 (.Y(N3144),.A(N651),.B(N2626));
AND2X1 AND2_691 (.Y(N3149),.A(N644),.B(N2619));
AND2X1 AND2_692 (.Y(N3155),.A(N2533),.B(N2269));
OR2X1 OR2_693 (.Y(N3159),.A(N1174),.B(N2878));
INVX1 NOT1_694 (.Y(N3167),.A(N2778));
AND2X1 AND2_695 (.Y(N3168),.A(N609),.B(N2508));
AND2X1 AND2_696 (.Y(N3169),.A(N604),.B(N2502));
AND2X1 AND2_697 (.Y(N3173),.A(N742),.B(N2496));
AND2X1 AND2_698 (.Y(N3178),.A(N734),.B(N2488));
AND2X1 AND2_699 (.Y(N3184),.A(N599),.B(N2482));
AND2X1 AND2_700 (.Y(N3185),.A(N727),.B(N2573));
AND2X1 AND2_701 (.Y(N3189),.A(N721),.B(N2567));
AND2X1 AND2_702 (.Y(N3195),.A(N715),.B(N2561));
AND2X1 AND2_703 (.Y(N3202),.A(N708),.B(N2554));
AND2X1 AND2_704 (.Y(N3210),.A(N609),.B(N2508));
AND2X1 AND2_705 (.Y(N3211),.A(N604),.B(N2502));
AND2X1 AND2_706 (.Y(N3215),.A(N742),.B(N2496));
AND2X1 AND2_707 (.Y(N3221),.A(N2488),.B(N734));
AND2X1 AND2_708 (.Y(N3228),.A(N599),.B(N2482));
AND2X1 AND2_709 (.Y(N3229),.A(N727),.B(N2573));
AND2X1 AND2_710 (.Y(N3232),.A(N721),.B(N2567));
AND2X1 AND2_711 (.Y(N3236),.A(N715),.B(N2561));
AND2X1 AND2_712 (.Y(N3241),.A(N708),.B(N2554));
OR2X1 OR2_713 (.Y(N3247),.A(N2913),.B(N2299));
OR2X1 OR2_714 (.Y(N3251),.A(N2914),.B(N2300));
OR2X1 OR2_715 (.Y(N3255),.A(N2915),.B(N2301));
OR2X1 OR2_716 (.Y(N3259),.A(N2916),.B(N2302));
OR2X1 OR2_717 (.Y(N3263),.A(N2917),.B(N2303));
OR2X1 OR2_718 (.Y(N3267),.A(N2918),.B(N2304));
OR2X1 OR2_719 (.Y(N3273),.A(N2919),.B(N2305));
OR2X1 OR2_720 (.Y(N3281),.A(N2920),.B(N2306));
OR2X1 OR2_721 (.Y(N3287),.A(N2921),.B(N2307));
OR2X1 OR2_722 (.Y(N3293),.A(N2922),.B(N2308));
OR2X1 OR2_723 (.Y(N3299),.A(N2924),.B(N2322));
OR2X1 OR2_724 (.Y(N3303),.A(N2925),.B(N2323));
OR2X1 OR2_725 (.Y(N3307),.A(N2926),.B(N2324));
OR2X1 OR2_726 (.Y(N3311),.A(N2927),.B(N2325));
OR2X1 OR2_727 (.Y(N3315),.A(N2929),.B(N2327));
OR2X1 OR2_728 (.Y(N3322),.A(N2930),.B(N2328));
OR2X1 OR2_729 (.Y(N3328),.A(N2931),.B(N2329));
OR2X1 OR2_730 (.Y(N3334),.A(N2932),.B(N2330));
OR2X1 OR2_731 (.Y(N3340),.A(N2934),.B(N2343));
OR2X1 OR2_732 (.Y(N3343),.A(N2935),.B(N2344));
OR2X1 OR2_733 (.Y(N3349),.A(N2936),.B(N2345));
OR2X1 OR2_734 (.Y(N3355),.A(N2937),.B(N2346));
AND2X1 AND2_735 (.Y(N3361),.A(N2761),.B(N2478));
AND2X1 AND2_736 (.Y(N3362),.A(N2757),.B(N2474));
AND2X1 AND2_737 (.Y(N3363),.A(N2753),.B(N2470));
AND2X1 AND2_738 (.Y(N3364),.A(N2749),.B(N2466));
AND2X1 AND2_739 (.Y(N3365),.A(N2745),.B(N2462));
AND2X1 AND2_740 (.Y(N3366),.A(N2741),.B(N2550));
AND2X1 AND2_741 (.Y(N3367),.A(N2737),.B(N2546));
AND2X1 AND2_742 (.Y(N3368),.A(N2733),.B(N2542));
AND2X1 AND2_743 (.Y(N3369),.A(N2729),.B(N2538));
AND2X1 AND2_744 (.Y(N3370),.A(N2670),.B(N2458));
AND2X1 AND2_745 (.Y(N3371),.A(N2666),.B(N2454));
AND2X1 AND2_746 (.Y(N3372),.A(N2662),.B(N2450));
AND2X1 AND2_747 (.Y(N3373),.A(N2658),.B(N2446));
AND2X1 AND2_748 (.Y(N3374),.A(N2654),.B(N2442));
AND2X1 AND2_749 (.Y(N3375),.A(N2988),.B(N2650));
AND2X1 AND2_750 (.Y(N3379),.A(N2650),.B(N1966));
INVX1 NOT1_751 (.Y(N3380),.A(N2781));
AND2X1 AND2_752 (.Y(N3381),.A(N695),.B(N2604));
OR2X1 OR2_753 (.Y(N3384),.A(N3005),.B(N2379));
OR2X1 OR2_754 (.Y(N3390),.A(N3006),.B(N2380));
OR2X1 OR2_755 (.Y(N3398),.A(N3007),.B(N2381));
OR2X1 OR2_756 (.Y(N3404),.A(N3008),.B(N2382));
OR2X1 OR2_757 (.Y(N3410),.A(N3009),.B(N2383));
OR2X1 OR2_758 (.Y(N3416),.A(N3021),.B(N2397));
OR2X1 OR2_759 (.Y(N3420),.A(N3022),.B(N2398));
OR2X1 OR2_760 (.Y(N3424),.A(N3023),.B(N2399));
OR2X1 OR2_761 (.Y(N3428),.A(N3024),.B(N2400));
OR2X1 OR2_762 (.Y(N3432),.A(N3025),.B(N2401));
OR2X1 OR2_763 (.Y(N3436),.A(N3026),.B(N2402));
OR2X1 OR2_764 (.Y(N3440),.A(N3027),.B(N2403));
OR2X1 OR2_765 (.Y(N3444),.A(N3028),.B(N2404));
OR2X1 OR2_766 (.Y(N3448),.A(N3029),.B(N2405));
INVX1 NOT1_767 (.Y(N3452),.A(N2790));
INVX1 NOT1_768 (.Y(N3453),.A(N2793));
OR2X1 OR2_769 (.Y(N3454),.A(N3034),.B(N2420));
OR2X1 OR2_770 (.Y(N3458),.A(N3035),.B(N2421));
OR2X1 OR2_771 (.Y(N3462),.A(N3036),.B(N2422));
OR2X1 OR2_772 (.Y(N3466),.A(N3037),.B(N2423));
OR2X1 OR2_773 (.Y(N3470),.A(N3038),.B(N2424));
OR2X1 OR2_774 (.Y(N3474),.A(N3039),.B(N2425));
OR2X1 OR2_775 (.Y(N3478),.A(N3040),.B(N2426));
OR2X1 OR2_776 (.Y(N3482),.A(N3041),.B(N2427));
INVX1 NOT1_777 (.Y(N3486),.A(N2796));
BUFX1 BUFF1_778 (.Y(N3487),.A(N2644));
BUFX1 BUFF1_779 (.Y(N3490),.A(N2638));
BUFX1 BUFF1_780 (.Y(N3493),.A(N2632));
BUFX1 BUFF1_781 (.Y(N3496),.A(N2626));
BUFX1 BUFF1_782 (.Y(N3499),.A(N2619));
BUFX1 BUFF1_783 (.Y(N3502),.A(N2523));
NOR2X1 NOR2_784 (.Y(N3507),.A(N1167),.B(N2868));
BUFX1 BUFF1_785 (.Y(N3510),.A(N2523));
NOR2X1 NOR2_786 (.Y(N3515),.A(N644),.B(N2619));
BUFX1 BUFF1_787 (.Y(N3518),.A(N2644));
BUFX1 BUFF1_788 (.Y(N3521),.A(N2638));
BUFX1 BUFF1_789 (.Y(N3524),.A(N2632));
BUFX1 BUFF1_790 (.Y(N3527),.A(N2626));
BUFX1 BUFF1_791 (.Y(N3530),.A(N2619));
BUFX1 BUFF1_792 (.Y(N3535),.A(N2619));
BUFX1 BUFF1_793 (.Y(N3539),.A(N2632));
BUFX1 BUFF1_794 (.Y(N3542),.A(N2626));
BUFX1 BUFF1_795 (.Y(N3545),.A(N2644));
BUFX1 BUFF1_796 (.Y(N3548),.A(N2638));
INVX1 NOT1_797 (.Y(N3551),.A(N2766));
INVX1 NOT1_798 (.Y(N3552),.A(N2769));
BUFX1 BUFF1_799 (.Y(N3553),.A(N2442));
BUFX1 BUFF1_800 (.Y(N3557),.A(N2450));
BUFX1 BUFF1_801 (.Y(N3560),.A(N2446));
BUFX1 BUFF1_802 (.Y(N3563),.A(N2458));
BUFX1 BUFF1_803 (.Y(N3566),.A(N2454));
INVX1 NOT1_804 (.Y(N3569),.A(N2772));
INVX1 NOT1_805 (.Y(N3570),.A(N2775));
BUFX1 BUFF1_806 (.Y(N3571),.A(N2554));
BUFX1 BUFF1_807 (.Y(N3574),.A(N2567));
BUFX1 BUFF1_808 (.Y(N3577),.A(N2561));
BUFX1 BUFF1_809 (.Y(N3580),.A(N2482));
BUFX1 BUFF1_810 (.Y(N3583),.A(N2573));
BUFX1 BUFF1_811 (.Y(N3586),.A(N2496));
BUFX1 BUFF1_812 (.Y(N3589),.A(N2488));
BUFX1 BUFF1_813 (.Y(N3592),.A(N2508));
BUFX1 BUFF1_814 (.Y(N3595),.A(N2502));
BUFX1 BUFF1_815 (.Y(N3598),.A(N2508));
BUFX1 BUFF1_816 (.Y(N3601),.A(N2502));
BUFX1 BUFF1_817 (.Y(N3604),.A(N2496));
BUFX1 BUFF1_818 (.Y(N3607),.A(N2482));
BUFX1 BUFF1_819 (.Y(N3610),.A(N2573));
BUFX1 BUFF1_820 (.Y(N3613),.A(N2567));
BUFX1 BUFF1_821 (.Y(N3616),.A(N2561));
BUFX1 BUFF1_822 (.Y(N3619),.A(N2488));
BUFX1 BUFF1_823 (.Y(N3622),.A(N2554));
NOR2X1 NOR2_824 (.Y(N3625),.A(N734),.B(N2488));
NOR2X1 NOR2_825 (.Y(N3628),.A(N708),.B(N2554));
BUFX1 BUFF1_826 (.Y(N3631),.A(N2508));
BUFX1 BUFF1_827 (.Y(N3634),.A(N2502));
BUFX1 BUFF1_828 (.Y(N3637),.A(N2496));
BUFX1 BUFF1_829 (.Y(N3640),.A(N2488));
BUFX1 BUFF1_830 (.Y(N3643),.A(N2482));
BUFX1 BUFF1_831 (.Y(N3646),.A(N2573));
BUFX1 BUFF1_832 (.Y(N3649),.A(N2567));
BUFX1 BUFF1_833 (.Y(N3652),.A(N2561));
BUFX1 BUFF1_834 (.Y(N3655),.A(N2554));
NOR2X1 NOR2_835 (.Y(N3658),.A(N2488),.B(N734));
BUFX1 BUFF1_836 (.Y(N3661),.A(N2674));
BUFX1 BUFF1_837 (.Y(N3664),.A(N2674));
BUFX1 BUFF1_838 (.Y(N3667),.A(N2761));
BUFX1 BUFF1_839 (.Y(N3670),.A(N2478));
BUFX1 BUFF1_840 (.Y(N3673),.A(N2757));
BUFX1 BUFF1_841 (.Y(N3676),.A(N2474));
BUFX1 BUFF1_842 (.Y(N3679),.A(N2753));
BUFX1 BUFF1_843 (.Y(N3682),.A(N2470));
BUFX1 BUFF1_844 (.Y(N3685),.A(N2745));
BUFX1 BUFF1_845 (.Y(N3688),.A(N2462));
BUFX1 BUFF1_846 (.Y(N3691),.A(N2741));
BUFX1 BUFF1_847 (.Y(N3694),.A(N2550));
BUFX1 BUFF1_848 (.Y(N3697),.A(N2737));
BUFX1 BUFF1_849 (.Y(N3700),.A(N2546));
BUFX1 BUFF1_850 (.Y(N3703),.A(N2733));
BUFX1 BUFF1_851 (.Y(N3706),.A(N2542));
BUFX1 BUFF1_852 (.Y(N3709),.A(N2749));
BUFX1 BUFF1_853 (.Y(N3712),.A(N2466));
BUFX1 BUFF1_854 (.Y(N3715),.A(N2729));
BUFX1 BUFF1_855 (.Y(N3718),.A(N2538));
BUFX1 BUFF1_856 (.Y(N3721),.A(N2704));
BUFX1 BUFF1_857 (.Y(N3724),.A(N2700));
BUFX1 BUFF1_858 (.Y(N3727),.A(N2696));
BUFX1 BUFF1_859 (.Y(N3730),.A(N2688));
BUFX1 BUFF1_860 (.Y(N3733),.A(N2692));
BUFX1 BUFF1_861 (.Y(N3736),.A(N2670));
BUFX1 BUFF1_862 (.Y(N3739),.A(N2458));
BUFX1 BUFF1_863 (.Y(N3742),.A(N2666));
BUFX1 BUFF1_864 (.Y(N3745),.A(N2454));
BUFX1 BUFF1_865 (.Y(N3748),.A(N2662));
BUFX1 BUFF1_866 (.Y(N3751),.A(N2450));
BUFX1 BUFF1_867 (.Y(N3754),.A(N2658));
BUFX1 BUFF1_868 (.Y(N3757),.A(N2446));
BUFX1 BUFF1_869 (.Y(N3760),.A(N2654));
BUFX1 BUFF1_870 (.Y(N3763),.A(N2442));
BUFX1 BUFF1_871 (.Y(N3766),.A(N2654));
BUFX1 BUFF1_872 (.Y(N3769),.A(N2662));
BUFX1 BUFF1_873 (.Y(N3772),.A(N2658));
BUFX1 BUFF1_874 (.Y(N3775),.A(N2670));
BUFX1 BUFF1_875 (.Y(N3778),.A(N2666));
INVX1 NOT1_876 (.Y(N3781),.A(N2784));
INVX1 NOT1_877 (.Y(N3782),.A(N2787));
OR2X1 OR2_878 (.Y(N3783),.A(N2928),.B(N2326));
OR2X1 OR2_879 (.Y(N3786),.A(N2933),.B(N2342));
OR2X1 OR2_880 (.Y(N3789),.A(N2923),.B(N2321));
BUFX1 BUFF1_881 (.Y(N3792),.A(N2688));
BUFX1 BUFF1_882 (.Y(N3795),.A(N2696));
BUFX1 BUFF1_883 (.Y(N3798),.A(N2692));
BUFX1 BUFF1_884 (.Y(N3801),.A(N2704));
BUFX1 BUFF1_885 (.Y(N3804),.A(N2700));
BUFX1 BUFF1_886 (.Y(N3807),.A(N2604));
BUFX1 BUFF1_887 (.Y(N3810),.A(N2611));
BUFX1 BUFF1_888 (.Y(N3813),.A(N2607));
BUFX1 BUFF1_889 (.Y(N3816),.A(N2615));
BUFX1 BUFF1_890 (.Y(N3819),.A(N2538));
BUFX1 BUFF1_891 (.Y(N3822),.A(N2546));
BUFX1 BUFF1_892 (.Y(N3825),.A(N2542));
BUFX1 BUFF1_893 (.Y(N3828),.A(N2462));
BUFX1 BUFF1_894 (.Y(N3831),.A(N2550));
BUFX1 BUFF1_895 (.Y(N3834),.A(N2470));
BUFX1 BUFF1_896 (.Y(N3837),.A(N2466));
BUFX1 BUFF1_897 (.Y(N3840),.A(N2478));
BUFX1 BUFF1_898 (.Y(N3843),.A(N2474));
BUFX1 BUFF1_899 (.Y(N3846),.A(N2615));
BUFX1 BUFF1_900 (.Y(N3849),.A(N2611));
BUFX1 BUFF1_901 (.Y(N3852),.A(N2607));
BUFX1 BUFF1_902 (.Y(N3855),.A(N2680));
BUFX1 BUFF1_903 (.Y(N3858),.A(N2729));
BUFX1 BUFF1_904 (.Y(N3861),.A(N2737));
BUFX1 BUFF1_905 (.Y(N3864),.A(N2733));
BUFX1 BUFF1_906 (.Y(N3867),.A(N2745));
BUFX1 BUFF1_907 (.Y(N3870),.A(N2741));
BUFX1 BUFF1_908 (.Y(N3873),.A(N2753));
BUFX1 BUFF1_909 (.Y(N3876),.A(N2749));
BUFX1 BUFF1_910 (.Y(N3879),.A(N2761));
BUFX1 BUFF1_911 (.Y(N3882),.A(N2757));
OR2X1 OR2_912 (.Y(N3885),.A(N3033),.B(N2419));
OR2X1 OR2_913 (.Y(N3888),.A(N3032),.B(N2418));
OR2X1 OR2_914 (.Y(N3891),.A(N3020),.B(N2396));
NAND2X1 NAND2_915 (.Y(N3953),.A(N3067),.B(N2117));
INVX1 NOT1_916 (.Y(N3954),.A(N3067));
NAND2X1 NAND2_917 (.Y(N3955),.A(N3070),.B(N2537));
INVX1 NOT1_918 (.Y(N3956),.A(N3070));
INVX1 NOT1_919 (.Y(N3958),.A(N3073));
INVX1 NOT1_920 (.Y(N3964),.A(N3080));
OR2X1 OR2_921 (.Y(N4193),.A(N1649),.B(N3379));
OR2X1 OR_tmp13 (.Y(ttmp13),.A(N2867),.B(N3130));
OR2X1 OR_tmp14 (.Y(N4303),.A(N1167),.B(ttmp13));
INVX1 NOT1_923 (.Y(N4308),.A(N3061));
INVX1 NOT1_924 (.Y(N4313),.A(N3064));
NAND2X1 NAND2_925 (.Y(N4326),.A(N2769),.B(N3551));
NAND2X1 NAND2_926 (.Y(N4327),.A(N2766),.B(N3552));
NAND2X1 NAND2_927 (.Y(N4333),.A(N2775),.B(N3569));
NAND2X1 NAND2_928 (.Y(N4334),.A(N2772),.B(N3570));
NAND2X1 NAND2_929 (.Y(N4411),.A(N2787),.B(N3781));
NAND2X1 NAND2_930 (.Y(N4412),.A(N2784),.B(N3782));
NAND2X1 NAND2_931 (.Y(N4463),.A(N3487),.B(N1828));
INVX1 NOT1_932 (.Y(N4464),.A(N3487));
NAND2X1 NAND2_933 (.Y(N4465),.A(N3490),.B(N1829));
INVX1 NOT1_934 (.Y(N4466),.A(N3490));
NAND2X1 NAND2_935 (.Y(N4467),.A(N3493),.B(N2267));
INVX1 NOT1_936 (.Y(N4468),.A(N3493));
NAND2X1 NAND2_937 (.Y(N4469),.A(N3496),.B(N1830));
INVX1 NOT1_938 (.Y(N4470),.A(N3496));
NAND2X1 NAND2_939 (.Y(N4471),.A(N3499),.B(N1833));
INVX1 NOT1_940 (.Y(N4472),.A(N3499));
INVX1 NOT1_941 (.Y(N4473),.A(N3122));
INVX1 NOT1_942 (.Y(N4474),.A(N3126));
NAND2X1 NAND2_943 (.Y(N4475),.A(N3518),.B(N1840));
INVX1 NOT1_944 (.Y(N4476),.A(N3518));
NAND2X1 NAND2_945 (.Y(N4477),.A(N3521),.B(N1841));
INVX1 NOT1_946 (.Y(N4478),.A(N3521));
NAND2X1 NAND2_947 (.Y(N4479),.A(N3524),.B(N2275));
INVX1 NOT1_948 (.Y(N4480),.A(N3524));
NAND2X1 NAND2_949 (.Y(N4481),.A(N3527),.B(N1842));
INVX1 NOT1_950 (.Y(N4482),.A(N3527));
NAND2X1 NAND2_951 (.Y(N4483),.A(N3530),.B(N1843));
INVX1 NOT1_952 (.Y(N4484),.A(N3530));
INVX1 NOT1_953 (.Y(N4485),.A(N3155));
INVX1 NOT1_954 (.Y(N4486),.A(N3159));
NAND2X1 NAND2_955 (.Y(N4487),.A(N1721),.B(N3954));
NAND2X1 NAND2_956 (.Y(N4488),.A(N2235),.B(N3956));
INVX1 NOT1_957 (.Y(N4489),.A(N3535));
NAND2X1 NAND2_958 (.Y(N4490),.A(N3535),.B(N3958));
INVX1 NOT1_959 (.Y(N4491),.A(N3539));
INVX1 NOT1_960 (.Y(N4492),.A(N3542));
INVX1 NOT1_961 (.Y(N4493),.A(N3545));
INVX1 NOT1_962 (.Y(N4494),.A(N3548));
INVX1 NOT1_963 (.Y(N4495),.A(N3553));
NAND2X1 NAND2_964 (.Y(N4496),.A(N3553),.B(N3964));
INVX1 NOT1_965 (.Y(N4497),.A(N3557));
INVX1 NOT1_966 (.Y(N4498),.A(N3560));
INVX1 NOT1_967 (.Y(N4499),.A(N3563));
INVX1 NOT1_968 (.Y(N4500),.A(N3566));
INVX1 NOT1_969 (.Y(N4501),.A(N3571));
NAND2X1 NAND2_970 (.Y(N4502),.A(N3571),.B(N3167));
INVX1 NOT1_971 (.Y(N4503),.A(N3574));
INVX1 NOT1_972 (.Y(N4504),.A(N3577));
INVX1 NOT1_973 (.Y(N4505),.A(N3580));
INVX1 NOT1_974 (.Y(N4506),.A(N3583));
NAND2X1 NAND2_975 (.Y(N4507),.A(N3598),.B(N1867));
INVX1 NOT1_976 (.Y(N4508),.A(N3598));
NAND2X1 NAND2_977 (.Y(N4509),.A(N3601),.B(N1868));
INVX1 NOT1_978 (.Y(N4510),.A(N3601));
NAND2X1 NAND2_979 (.Y(N4511),.A(N3604),.B(N1869));
INVX1 NOT1_980 (.Y(N4512),.A(N3604));
NAND2X1 NAND2_981 (.Y(N4513),.A(N3607),.B(N1870));
INVX1 NOT1_982 (.Y(N4514),.A(N3607));
NAND2X1 NAND2_983 (.Y(N4515),.A(N3610),.B(N1871));
INVX1 NOT1_984 (.Y(N4516),.A(N3610));
NAND2X1 NAND2_985 (.Y(N4517),.A(N3613),.B(N1872));
INVX1 NOT1_986 (.Y(N4518),.A(N3613));
NAND2X1 NAND2_987 (.Y(N4519),.A(N3616),.B(N1873));
INVX1 NOT1_988 (.Y(N4520),.A(N3616));
NAND2X1 NAND2_989 (.Y(N4521),.A(N3619),.B(N1874));
INVX1 NOT1_990 (.Y(N4522),.A(N3619));
NAND2X1 NAND2_991 (.Y(N4523),.A(N3622),.B(N1875));
INVX1 NOT1_992 (.Y(N4524),.A(N3622));
NAND2X1 NAND2_993 (.Y(N4525),.A(N3631),.B(N1876));
INVX1 NOT1_994 (.Y(N4526),.A(N3631));
NAND2X1 NAND2_995 (.Y(N4527),.A(N3634),.B(N1877));
INVX1 NOT1_996 (.Y(N4528),.A(N3634));
NAND2X1 NAND2_997 (.Y(N4529),.A(N3637),.B(N1878));
INVX1 NOT1_998 (.Y(N4530),.A(N3637));
NAND2X1 NAND2_999 (.Y(N4531),.A(N3640),.B(N1879));
INVX1 NOT1_1000 (.Y(N4532),.A(N3640));
NAND2X1 NAND2_1001 (.Y(N4533),.A(N3643),.B(N1880));
INVX1 NOT1_1002 (.Y(N4534),.A(N3643));
NAND2X1 NAND2_1003 (.Y(N4535),.A(N3646),.B(N1881));
INVX1 NOT1_1004 (.Y(N4536),.A(N3646));
NAND2X1 NAND2_1005 (.Y(N4537),.A(N3649),.B(N1882));
INVX1 NOT1_1006 (.Y(N4538),.A(N3649));
NAND2X1 NAND2_1007 (.Y(N4539),.A(N3652),.B(N1883));
INVX1 NOT1_1008 (.Y(N4540),.A(N3652));
NAND2X1 NAND2_1009 (.Y(N4541),.A(N3655),.B(N1884));
INVX1 NOT1_1010 (.Y(N4542),.A(N3655));
INVX1 NOT1_1011 (.Y(N4543),.A(N3658));
AND2X1 AND2_1012 (.Y(N4544),.A(N806),.B(N3293));
AND2X1 AND2_1013 (.Y(N4545),.A(N800),.B(N3287));
AND2X1 AND2_1014 (.Y(N4549),.A(N794),.B(N3281));
AND2X1 AND2_1015 (.Y(N4555),.A(N3273),.B(N786));
AND2X1 AND2_1016 (.Y(N4562),.A(N780),.B(N3267));
AND2X1 AND2_1017 (.Y(N4563),.A(N774),.B(N3355));
AND2X1 AND2_1018 (.Y(N4566),.A(N768),.B(N3349));
AND2X1 AND2_1019 (.Y(N4570),.A(N762),.B(N3343));
INVX1 NOT1_1020 (.Y(N4575),.A(N3661));
AND2X1 AND2_1021 (.Y(N4576),.A(N806),.B(N3293));
AND2X1 AND2_1022 (.Y(N4577),.A(N800),.B(N3287));
AND2X1 AND2_1023 (.Y(N4581),.A(N794),.B(N3281));
AND2X1 AND2_1024 (.Y(N4586),.A(N786),.B(N3273));
AND2X1 AND2_1025 (.Y(N4592),.A(N780),.B(N3267));
AND2X1 AND2_1026 (.Y(N4593),.A(N774),.B(N3355));
AND2X1 AND2_1027 (.Y(N4597),.A(N768),.B(N3349));
AND2X1 AND2_1028 (.Y(N4603),.A(N762),.B(N3343));
INVX1 NOT1_1029 (.Y(N4610),.A(N3664));
INVX1 NOT1_1030 (.Y(N4611),.A(N3667));
INVX1 NOT1_1031 (.Y(N4612),.A(N3670));
INVX1 NOT1_1032 (.Y(N4613),.A(N3673));
INVX1 NOT1_1033 (.Y(N4614),.A(N3676));
INVX1 NOT1_1034 (.Y(N4615),.A(N3679));
INVX1 NOT1_1035 (.Y(N4616),.A(N3682));
INVX1 NOT1_1036 (.Y(N4617),.A(N3685));
INVX1 NOT1_1037 (.Y(N4618),.A(N3688));
INVX1 NOT1_1038 (.Y(N4619),.A(N3691));
INVX1 NOT1_1039 (.Y(N4620),.A(N3694));
INVX1 NOT1_1040 (.Y(N4621),.A(N3697));
INVX1 NOT1_1041 (.Y(N4622),.A(N3700));
INVX1 NOT1_1042 (.Y(N4623),.A(N3703));
INVX1 NOT1_1043 (.Y(N4624),.A(N3706));
INVX1 NOT1_1044 (.Y(N4625),.A(N3709));
INVX1 NOT1_1045 (.Y(N4626),.A(N3712));
INVX1 NOT1_1046 (.Y(N4627),.A(N3715));
INVX1 NOT1_1047 (.Y(N4628),.A(N3718));
INVX1 NOT1_1048 (.Y(N4629),.A(N3721));
AND2X1 AND2_1049 (.Y(N4630),.A(N3448),.B(N2704));
INVX1 NOT1_1050 (.Y(N4631),.A(N3724));
AND2X1 AND2_1051 (.Y(N4632),.A(N3444),.B(N2700));
INVX1 NOT1_1052 (.Y(N4633),.A(N3727));
AND2X1 AND2_1053 (.Y(N4634),.A(N3440),.B(N2696));
AND2X1 AND2_1054 (.Y(N4635),.A(N3436),.B(N2692));
INVX1 NOT1_1055 (.Y(N4636),.A(N3730));
AND2X1 AND2_1056 (.Y(N4637),.A(N3432),.B(N2688));
AND2X1 AND2_1057 (.Y(N4638),.A(N3428),.B(N3311));
AND2X1 AND2_1058 (.Y(N4639),.A(N3424),.B(N3307));
AND2X1 AND2_1059 (.Y(N4640),.A(N3420),.B(N3303));
AND2X1 AND2_1060 (.Y(N4641),.A(N3416),.B(N3299));
INVX1 NOT1_1061 (.Y(N4642),.A(N3733));
INVX1 NOT1_1062 (.Y(N4643),.A(N3736));
INVX1 NOT1_1063 (.Y(N4644),.A(N3739));
INVX1 NOT1_1064 (.Y(N4645),.A(N3742));
INVX1 NOT1_1065 (.Y(N4646),.A(N3745));
INVX1 NOT1_1066 (.Y(N4647),.A(N3748));
INVX1 NOT1_1067 (.Y(N4648),.A(N3751));
INVX1 NOT1_1068 (.Y(N4649),.A(N3754));
INVX1 NOT1_1069 (.Y(N4650),.A(N3757));
INVX1 NOT1_1070 (.Y(N4651),.A(N3760));
INVX1 NOT1_1071 (.Y(N4652),.A(N3763));
INVX1 NOT1_1072 (.Y(N4653),.A(N3375));
AND2X1 AND2_1073 (.Y(N4656),.A(N865),.B(N3410));
AND2X1 AND2_1074 (.Y(N4657),.A(N859),.B(N3404));
AND2X1 AND2_1075 (.Y(N4661),.A(N853),.B(N3398));
AND2X1 AND2_1076 (.Y(N4667),.A(N3390),.B(N845));
AND2X1 AND2_1077 (.Y(N4674),.A(N839),.B(N3384));
AND2X1 AND2_1078 (.Y(N4675),.A(N833),.B(N3334));
AND2X1 AND2_1079 (.Y(N4678),.A(N827),.B(N3328));
AND2X1 AND2_1080 (.Y(N4682),.A(N821),.B(N3322));
AND2X1 AND2_1081 (.Y(N4687),.A(N814),.B(N3315));
INVX1 NOT1_1082 (.Y(N4693),.A(N3766));
NAND2X1 NAND2_1083 (.Y(N4694),.A(N3766),.B(N3380));
INVX1 NOT1_1084 (.Y(N4695),.A(N3769));
INVX1 NOT1_1085 (.Y(N4696),.A(N3772));
INVX1 NOT1_1086 (.Y(N4697),.A(N3775));
INVX1 NOT1_1087 (.Y(N4698),.A(N3778));
INVX1 NOT1_1088 (.Y(N4699),.A(N3783));
INVX1 NOT1_1089 (.Y(N4700),.A(N3786));
AND2X1 AND2_1090 (.Y(N4701),.A(N865),.B(N3410));
AND2X1 AND2_1091 (.Y(N4702),.A(N859),.B(N3404));
AND2X1 AND2_1092 (.Y(N4706),.A(N853),.B(N3398));
AND2X1 AND2_1093 (.Y(N4711),.A(N845),.B(N3390));
AND2X1 AND2_1094 (.Y(N4717),.A(N839),.B(N3384));
AND2X1 AND2_1095 (.Y(N4718),.A(N833),.B(N3334));
AND2X1 AND2_1096 (.Y(N4722),.A(N827),.B(N3328));
AND2X1 AND2_1097 (.Y(N4728),.A(N821),.B(N3322));
AND2X1 AND2_1098 (.Y(N4735),.A(N814),.B(N3315));
INVX1 NOT1_1099 (.Y(N4743),.A(N3789));
INVX1 NOT1_1100 (.Y(N4744),.A(N3792));
INVX1 NOT1_1101 (.Y(N4745),.A(N3807));
NAND2X1 NAND2_1102 (.Y(N4746),.A(N3807),.B(N3452));
INVX1 NOT1_1103 (.Y(N4747),.A(N3810));
INVX1 NOT1_1104 (.Y(N4748),.A(N3813));
INVX1 NOT1_1105 (.Y(N4749),.A(N3816));
INVX1 NOT1_1106 (.Y(N4750),.A(N3819));
NAND2X1 NAND2_1107 (.Y(N4751),.A(N3819),.B(N3453));
INVX1 NOT1_1108 (.Y(N4752),.A(N3822));
INVX1 NOT1_1109 (.Y(N4753),.A(N3825));
INVX1 NOT1_1110 (.Y(N4754),.A(N3828));
INVX1 NOT1_1111 (.Y(N4755),.A(N3831));
AND2X1 AND2_1112 (.Y(N4756),.A(N3482),.B(N3263));
AND2X1 AND2_1113 (.Y(N4757),.A(N3478),.B(N3259));
AND2X1 AND2_1114 (.Y(N4758),.A(N3474),.B(N3255));
AND2X1 AND2_1115 (.Y(N4759),.A(N3470),.B(N3251));
AND2X1 AND2_1116 (.Y(N4760),.A(N3466),.B(N3247));
INVX1 NOT1_1117 (.Y(N4761),.A(N3846));
AND2X1 AND2_1118 (.Y(N4762),.A(N3462),.B(N2615));
INVX1 NOT1_1119 (.Y(N4763),.A(N3849));
AND2X1 AND2_1120 (.Y(N4764),.A(N3458),.B(N2611));
INVX1 NOT1_1121 (.Y(N4765),.A(N3852));
AND2X1 AND2_1122 (.Y(N4766),.A(N3454),.B(N2607));
AND2X1 AND2_1123 (.Y(N4767),.A(N2680),.B(N3381));
INVX1 NOT1_1124 (.Y(N4768),.A(N3855));
AND2X1 AND2_1125 (.Y(N4769),.A(N3340),.B(N695));
INVX1 NOT1_1126 (.Y(N4775),.A(N3858));
NAND2X1 NAND2_1127 (.Y(N4776),.A(N3858),.B(N3486));
INVX1 NOT1_1128 (.Y(N4777),.A(N3861));
INVX1 NOT1_1129 (.Y(N4778),.A(N3864));
INVX1 NOT1_1130 (.Y(N4779),.A(N3867));
INVX1 NOT1_1131 (.Y(N4780),.A(N3870));
INVX1 NOT1_1132 (.Y(N4781),.A(N3885));
INVX1 NOT1_1133 (.Y(N4782),.A(N3888));
INVX1 NOT1_1134 (.Y(N4783),.A(N3891));
OR2X1 OR2_1135 (.Y(N4784),.A(N3131),.B(N3134));
INVX1 NOT1_1136 (.Y(N4789),.A(N3502));
INVX1 NOT1_1137 (.Y(N4790),.A(N3131));
INVX1 NOT1_1138 (.Y(N4793),.A(N3507));
INVX1 NOT1_1139 (.Y(N4794),.A(N3510));
INVX1 NOT1_1140 (.Y(N4795),.A(N3515));
BUFX1 BUFF1_1141 (.Y(N4796),.A(N3114));
INVX1 NOT1_1142 (.Y(N4799),.A(N3586));
INVX1 NOT1_1143 (.Y(N4800),.A(N3589));
INVX1 NOT1_1144 (.Y(N4801),.A(N3592));
INVX1 NOT1_1145 (.Y(N4802),.A(N3595));
NAND2X1 NAND2_1146 (.Y(N4803),.A(N4326),.B(N4327));
NAND2X1 NAND2_1147 (.Y(N4806),.A(N4333),.B(N4334));
INVX1 NOT1_1148 (.Y(N4809),.A(N3625));
BUFX1 BUFF1_1149 (.Y(N4810),.A(N3178));
INVX1 NOT1_1150 (.Y(N4813),.A(N3628));
BUFX1 BUFF1_1151 (.Y(N4814),.A(N3202));
BUFX1 BUFF1_1152 (.Y(N4817),.A(N3221));
BUFX1 BUFF1_1153 (.Y(N4820),.A(N3293));
BUFX1 BUFF1_1154 (.Y(N4823),.A(N3287));
BUFX1 BUFF1_1155 (.Y(N4826),.A(N3281));
BUFX1 BUFF1_1156 (.Y(N4829),.A(N3273));
BUFX1 BUFF1_1157 (.Y(N4832),.A(N3267));
BUFX1 BUFF1_1158 (.Y(N4835),.A(N3355));
BUFX1 BUFF1_1159 (.Y(N4838),.A(N3349));
BUFX1 BUFF1_1160 (.Y(N4841),.A(N3343));
NOR2X1 NOR2_1161 (.Y(N4844),.A(N3273),.B(N786));
BUFX1 BUFF1_1162 (.Y(N4847),.A(N3293));
BUFX1 BUFF1_1163 (.Y(N4850),.A(N3287));
BUFX1 BUFF1_1164 (.Y(N4853),.A(N3281));
BUFX1 BUFF1_1165 (.Y(N4856),.A(N3267));
BUFX1 BUFF1_1166 (.Y(N4859),.A(N3355));
BUFX1 BUFF1_1167 (.Y(N4862),.A(N3349));
BUFX1 BUFF1_1168 (.Y(N4865),.A(N3343));
BUFX1 BUFF1_1169 (.Y(N4868),.A(N3273));
NOR2X1 NOR2_1170 (.Y(N4871),.A(N786),.B(N3273));
BUFX1 BUFF1_1171 (.Y(N4874),.A(N3448));
BUFX1 BUFF1_1172 (.Y(N4877),.A(N3444));
BUFX1 BUFF1_1173 (.Y(N4880),.A(N3440));
BUFX1 BUFF1_1174 (.Y(N4883),.A(N3432));
BUFX1 BUFF1_1175 (.Y(N4886),.A(N3428));
BUFX1 BUFF1_1176 (.Y(N4889),.A(N3311));
BUFX1 BUFF1_1177 (.Y(N4892),.A(N3424));
BUFX1 BUFF1_1178 (.Y(N4895),.A(N3307));
BUFX1 BUFF1_1179 (.Y(N4898),.A(N3420));
BUFX1 BUFF1_1180 (.Y(N4901),.A(N3303));
BUFX1 BUFF1_1181 (.Y(N4904),.A(N3436));
BUFX1 BUFF1_1182 (.Y(N4907),.A(N3416));
BUFX1 BUFF1_1183 (.Y(N4910),.A(N3299));
BUFX1 BUFF1_1184 (.Y(N4913),.A(N3410));
BUFX1 BUFF1_1185 (.Y(N4916),.A(N3404));
BUFX1 BUFF1_1186 (.Y(N4919),.A(N3398));
BUFX1 BUFF1_1187 (.Y(N4922),.A(N3390));
BUFX1 BUFF1_1188 (.Y(N4925),.A(N3384));
BUFX1 BUFF1_1189 (.Y(N4928),.A(N3334));
BUFX1 BUFF1_1190 (.Y(N4931),.A(N3328));
BUFX1 BUFF1_1191 (.Y(N4934),.A(N3322));
BUFX1 BUFF1_1192 (.Y(N4937),.A(N3315));
NOR2X1 NOR2_1193 (.Y(N4940),.A(N3390),.B(N845));
BUFX1 BUFF1_1194 (.Y(N4943),.A(N3315));
BUFX1 BUFF1_1195 (.Y(N4946),.A(N3328));
BUFX1 BUFF1_1196 (.Y(N4949),.A(N3322));
BUFX1 BUFF1_1197 (.Y(N4952),.A(N3384));
BUFX1 BUFF1_1198 (.Y(N4955),.A(N3334));
BUFX1 BUFF1_1199 (.Y(N4958),.A(N3398));
BUFX1 BUFF1_1200 (.Y(N4961),.A(N3390));
BUFX1 BUFF1_1201 (.Y(N4964),.A(N3410));
BUFX1 BUFF1_1202 (.Y(N4967),.A(N3404));
BUFX1 BUFF1_1203 (.Y(N4970),.A(N3340));
BUFX1 BUFF1_1204 (.Y(N4973),.A(N3349));
BUFX1 BUFF1_1205 (.Y(N4976),.A(N3343));
BUFX1 BUFF1_1206 (.Y(N4979),.A(N3267));
BUFX1 BUFF1_1207 (.Y(N4982),.A(N3355));
BUFX1 BUFF1_1208 (.Y(N4985),.A(N3281));
BUFX1 BUFF1_1209 (.Y(N4988),.A(N3273));
BUFX1 BUFF1_1210 (.Y(N4991),.A(N3293));
BUFX1 BUFF1_1211 (.Y(N4994),.A(N3287));
NAND2X1 NAND2_1212 (.Y(N4997),.A(N4411),.B(N4412));
BUFX1 BUFF1_1213 (.Y(N5000),.A(N3410));
BUFX1 BUFF1_1214 (.Y(N5003),.A(N3404));
BUFX1 BUFF1_1215 (.Y(N5006),.A(N3398));
BUFX1 BUFF1_1216 (.Y(N5009),.A(N3384));
BUFX1 BUFF1_1217 (.Y(N5012),.A(N3334));
BUFX1 BUFF1_1218 (.Y(N5015),.A(N3328));
BUFX1 BUFF1_1219 (.Y(N5018),.A(N3322));
BUFX1 BUFF1_1220 (.Y(N5021),.A(N3390));
BUFX1 BUFF1_1221 (.Y(N5024),.A(N3315));
NOR2X1 NOR2_1222 (.Y(N5027),.A(N845),.B(N3390));
NOR2X1 NOR2_1223 (.Y(N5030),.A(N814),.B(N3315));
BUFX1 BUFF1_1224 (.Y(N5033),.A(N3299));
BUFX1 BUFF1_1225 (.Y(N5036),.A(N3307));
BUFX1 BUFF1_1226 (.Y(N5039),.A(N3303));
BUFX1 BUFF1_1227 (.Y(N5042),.A(N3311));
INVX1 NOT1_1228 (.Y(N5045),.A(N3795));
INVX1 NOT1_1229 (.Y(N5046),.A(N3798));
INVX1 NOT1_1230 (.Y(N5047),.A(N3801));
INVX1 NOT1_1231 (.Y(N5048),.A(N3804));
BUFX1 BUFF1_1232 (.Y(N5049),.A(N3247));
BUFX1 BUFF1_1233 (.Y(N5052),.A(N3255));
BUFX1 BUFF1_1234 (.Y(N5055),.A(N3251));
BUFX1 BUFF1_1235 (.Y(N5058),.A(N3263));
BUFX1 BUFF1_1236 (.Y(N5061),.A(N3259));
INVX1 NOT1_1237 (.Y(N5064),.A(N3834));
INVX1 NOT1_1238 (.Y(N5065),.A(N3837));
INVX1 NOT1_1239 (.Y(N5066),.A(N3840));
INVX1 NOT1_1240 (.Y(N5067),.A(N3843));
BUFX1 BUFF1_1241 (.Y(N5068),.A(N3482));
BUFX1 BUFF1_1242 (.Y(N5071),.A(N3263));
BUFX1 BUFF1_1243 (.Y(N5074),.A(N3478));
BUFX1 BUFF1_1244 (.Y(N5077),.A(N3259));
BUFX1 BUFF1_1245 (.Y(N5080),.A(N3474));
BUFX1 BUFF1_1246 (.Y(N5083),.A(N3255));
BUFX1 BUFF1_1247 (.Y(N5086),.A(N3466));
BUFX1 BUFF1_1248 (.Y(N5089),.A(N3247));
BUFX1 BUFF1_1249 (.Y(N5092),.A(N3462));
BUFX1 BUFF1_1250 (.Y(N5095),.A(N3458));
BUFX1 BUFF1_1251 (.Y(N5098),.A(N3454));
BUFX1 BUFF1_1252 (.Y(N5101),.A(N3470));
BUFX1 BUFF1_1253 (.Y(N5104),.A(N3251));
BUFX1 BUFF1_1254 (.Y(N5107),.A(N3381));
INVX1 NOT1_1255 (.Y(N5110),.A(N3873));
INVX1 NOT1_1256 (.Y(N5111),.A(N3876));
INVX1 NOT1_1257 (.Y(N5112),.A(N3879));
INVX1 NOT1_1258 (.Y(N5113),.A(N3882));
BUFX1 BUFF1_1259 (.Y(N5114),.A(N3458));
BUFX1 BUFF1_1260 (.Y(N5117),.A(N3454));
BUFX1 BUFF1_1261 (.Y(N5120),.A(N3466));
BUFX1 BUFF1_1262 (.Y(N5123),.A(N3462));
BUFX1 BUFF1_1263 (.Y(N5126),.A(N3474));
BUFX1 BUFF1_1264 (.Y(N5129),.A(N3470));
BUFX1 BUFF1_1265 (.Y(N5132),.A(N3482));
BUFX1 BUFF1_1266 (.Y(N5135),.A(N3478));
BUFX1 BUFF1_1267 (.Y(N5138),.A(N3416));
BUFX1 BUFF1_1268 (.Y(N5141),.A(N3424));
BUFX1 BUFF1_1269 (.Y(N5144),.A(N3420));
BUFX1 BUFF1_1270 (.Y(N5147),.A(N3432));
BUFX1 BUFF1_1271 (.Y(N5150),.A(N3428));
BUFX1 BUFF1_1272 (.Y(N5153),.A(N3440));
BUFX1 BUFF1_1273 (.Y(N5156),.A(N3436));
BUFX1 BUFF1_1274 (.Y(N5159),.A(N3448));
BUFX1 BUFF1_1275 (.Y(N5162),.A(N3444));
NAND2X1 NAND2_1276 (.Y(N5165),.A(N4486),.B(N4485));
NAND2X1 NAND2_1277 (.Y(N5166),.A(N4474),.B(N4473));
NAND2X1 NAND2_1278 (.Y(N5167),.A(N1290),.B(N4464));
NAND2X1 NAND2_1279 (.Y(N5168),.A(N1293),.B(N4466));
NAND2X1 NAND2_1280 (.Y(N5169),.A(N2074),.B(N4468));
NAND2X1 NAND2_1281 (.Y(N5170),.A(N1296),.B(N4470));
NAND2X1 NAND2_1282 (.Y(N5171),.A(N1302),.B(N4472));
NAND2X1 NAND2_1283 (.Y(N5172),.A(N1314),.B(N4476));
NAND2X1 NAND2_1284 (.Y(N5173),.A(N1317),.B(N4478));
NAND2X1 NAND2_1285 (.Y(N5174),.A(N2081),.B(N4480));
NAND2X1 NAND2_1286 (.Y(N5175),.A(N1320),.B(N4482));
NAND2X1 NAND2_1287 (.Y(N5176),.A(N1323),.B(N4484));
NAND2X1 NAND2_1288 (.Y(N5177),.A(N3953),.B(N4487));
NAND2X1 NAND2_1289 (.Y(N5178),.A(N3955),.B(N4488));
NAND2X1 NAND2_1290 (.Y(N5179),.A(N3073),.B(N4489));
NAND2X1 NAND2_1291 (.Y(N5180),.A(N3542),.B(N4491));
NAND2X1 NAND2_1292 (.Y(N5181),.A(N3539),.B(N4492));
NAND2X1 NAND2_1293 (.Y(N5182),.A(N3548),.B(N4493));
NAND2X1 NAND2_1294 (.Y(N5183),.A(N3545),.B(N4494));
NAND2X1 NAND2_1295 (.Y(N5184),.A(N3080),.B(N4495));
NAND2X1 NAND2_1296 (.Y(N5185),.A(N3560),.B(N4497));
NAND2X1 NAND2_1297 (.Y(N5186),.A(N3557),.B(N4498));
NAND2X1 NAND2_1298 (.Y(N5187),.A(N3566),.B(N4499));
NAND2X1 NAND2_1299 (.Y(N5188),.A(N3563),.B(N4500));
NAND2X1 NAND2_1300 (.Y(N5189),.A(N2778),.B(N4501));
NAND2X1 NAND2_1301 (.Y(N5190),.A(N3577),.B(N4503));
NAND2X1 NAND2_1302 (.Y(N5191),.A(N3574),.B(N4504));
NAND2X1 NAND2_1303 (.Y(N5192),.A(N3583),.B(N4505));
NAND2X1 NAND2_1304 (.Y(N5193),.A(N3580),.B(N4506));
NAND2X1 NAND2_1305 (.Y(N5196),.A(N1326),.B(N4508));
NAND2X1 NAND2_1306 (.Y(N5197),.A(N1329),.B(N4510));
NAND2X1 NAND2_1307 (.Y(N5198),.A(N1332),.B(N4512));
NAND2X1 NAND2_1308 (.Y(N5199),.A(N1335),.B(N4514));
NAND2X1 NAND2_1309 (.Y(N5200),.A(N1338),.B(N4516));
NAND2X1 NAND2_1310 (.Y(N5201),.A(N1341),.B(N4518));
NAND2X1 NAND2_1311 (.Y(N5202),.A(N1344),.B(N4520));
NAND2X1 NAND2_1312 (.Y(N5203),.A(N1347),.B(N4522));
NAND2X1 NAND2_1313 (.Y(N5204),.A(N1350),.B(N4524));
NAND2X1 NAND2_1314 (.Y(N5205),.A(N1353),.B(N4526));
NAND2X1 NAND2_1315 (.Y(N5206),.A(N1356),.B(N4528));
NAND2X1 NAND2_1316 (.Y(N5207),.A(N1359),.B(N4530));
NAND2X1 NAND2_1317 (.Y(N5208),.A(N1362),.B(N4532));
NAND2X1 NAND2_1318 (.Y(N5209),.A(N1365),.B(N4534));
NAND2X1 NAND2_1319 (.Y(N5210),.A(N1368),.B(N4536));
NAND2X1 NAND2_1320 (.Y(N5211),.A(N1371),.B(N4538));
NAND2X1 NAND2_1321 (.Y(N5212),.A(N1374),.B(N4540));
NAND2X1 NAND2_1322 (.Y(N5213),.A(N1377),.B(N4542));
NAND2X1 NAND2_1323 (.Y(N5283),.A(N3670),.B(N4611));
NAND2X1 NAND2_1324 (.Y(N5284),.A(N3667),.B(N4612));
NAND2X1 NAND2_1325 (.Y(N5285),.A(N3676),.B(N4613));
NAND2X1 NAND2_1326 (.Y(N5286),.A(N3673),.B(N4614));
NAND2X1 NAND2_1327 (.Y(N5287),.A(N3682),.B(N4615));
NAND2X1 NAND2_1328 (.Y(N5288),.A(N3679),.B(N4616));
NAND2X1 NAND2_1329 (.Y(N5289),.A(N3688),.B(N4617));
NAND2X1 NAND2_1330 (.Y(N5290),.A(N3685),.B(N4618));
NAND2X1 NAND2_1331 (.Y(N5291),.A(N3694),.B(N4619));
NAND2X1 NAND2_1332 (.Y(N5292),.A(N3691),.B(N4620));
NAND2X1 NAND2_1333 (.Y(N5293),.A(N3700),.B(N4621));
NAND2X1 NAND2_1334 (.Y(N5294),.A(N3697),.B(N4622));
NAND2X1 NAND2_1335 (.Y(N5295),.A(N3706),.B(N4623));
NAND2X1 NAND2_1336 (.Y(N5296),.A(N3703),.B(N4624));
NAND2X1 NAND2_1337 (.Y(N5297),.A(N3712),.B(N4625));
NAND2X1 NAND2_1338 (.Y(N5298),.A(N3709),.B(N4626));
NAND2X1 NAND2_1339 (.Y(N5299),.A(N3718),.B(N4627));
NAND2X1 NAND2_1340 (.Y(N5300),.A(N3715),.B(N4628));
NAND2X1 NAND2_1341 (.Y(N5314),.A(N3739),.B(N4643));
NAND2X1 NAND2_1342 (.Y(N5315),.A(N3736),.B(N4644));
NAND2X1 NAND2_1343 (.Y(N5316),.A(N3745),.B(N4645));
NAND2X1 NAND2_1344 (.Y(N5317),.A(N3742),.B(N4646));
NAND2X1 NAND2_1345 (.Y(N5318),.A(N3751),.B(N4647));
NAND2X1 NAND2_1346 (.Y(N5319),.A(N3748),.B(N4648));
NAND2X1 NAND2_1347 (.Y(N5320),.A(N3757),.B(N4649));
NAND2X1 NAND2_1348 (.Y(N5321),.A(N3754),.B(N4650));
NAND2X1 NAND2_1349 (.Y(N5322),.A(N3763),.B(N4651));
NAND2X1 NAND2_1350 (.Y(N5323),.A(N3760),.B(N4652));
INVX1 NOT1_1351 (.Y(N5324),.A(N4193));
NAND2X1 NAND2_1352 (.Y(N5363),.A(N2781),.B(N4693));
NAND2X1 NAND2_1353 (.Y(N5364),.A(N3772),.B(N4695));
NAND2X1 NAND2_1354 (.Y(N5365),.A(N3769),.B(N4696));
NAND2X1 NAND2_1355 (.Y(N5366),.A(N3778),.B(N4697));
NAND2X1 NAND2_1356 (.Y(N5367),.A(N3775),.B(N4698));
NAND2X1 NAND2_1357 (.Y(N5425),.A(N2790),.B(N4745));
NAND2X1 NAND2_1358 (.Y(N5426),.A(N3813),.B(N4747));
NAND2X1 NAND2_1359 (.Y(N5427),.A(N3810),.B(N4748));
NAND2X1 NAND2_1360 (.Y(N5429),.A(N2793),.B(N4750));
NAND2X1 NAND2_1361 (.Y(N5430),.A(N3825),.B(N4752));
NAND2X1 NAND2_1362 (.Y(N5431),.A(N3822),.B(N4753));
NAND2X1 NAND2_1363 (.Y(N5432),.A(N3831),.B(N4754));
NAND2X1 NAND2_1364 (.Y(N5433),.A(N3828),.B(N4755));
NAND2X1 NAND2_1365 (.Y(N5451),.A(N2796),.B(N4775));
NAND2X1 NAND2_1366 (.Y(N5452),.A(N3864),.B(N4777));
NAND2X1 NAND2_1367 (.Y(N5453),.A(N3861),.B(N4778));
NAND2X1 NAND2_1368 (.Y(N5454),.A(N3870),.B(N4779));
NAND2X1 NAND2_1369 (.Y(N5455),.A(N3867),.B(N4780));
NAND2X1 NAND2_1370 (.Y(N5456),.A(N3888),.B(N4781));
NAND2X1 NAND2_1371 (.Y(N5457),.A(N3885),.B(N4782));
INVX1 NOT1_1372 (.Y(N5469),.A(N4303));
NAND2X1 NAND2_1373 (.Y(N5474),.A(N3589),.B(N4799));
NAND2X1 NAND2_1374 (.Y(N5475),.A(N3586),.B(N4800));
NAND2X1 NAND2_1375 (.Y(N5476),.A(N3595),.B(N4801));
NAND2X1 NAND2_1376 (.Y(N5477),.A(N3592),.B(N4802));
NAND2X1 NAND2_1377 (.Y(N5571),.A(N3798),.B(N5045));
NAND2X1 NAND2_1378 (.Y(N5572),.A(N3795),.B(N5046));
NAND2X1 NAND2_1379 (.Y(N5573),.A(N3804),.B(N5047));
NAND2X1 NAND2_1380 (.Y(N5574),.A(N3801),.B(N5048));
NAND2X1 NAND2_1381 (.Y(N5584),.A(N3837),.B(N5064));
NAND2X1 NAND2_1382 (.Y(N5585),.A(N3834),.B(N5065));
NAND2X1 NAND2_1383 (.Y(N5586),.A(N3843),.B(N5066));
NAND2X1 NAND2_1384 (.Y(N5587),.A(N3840),.B(N5067));
NAND2X1 NAND2_1385 (.Y(N5602),.A(N3876),.B(N5110));
NAND2X1 NAND2_1386 (.Y(N5603),.A(N3873),.B(N5111));
NAND2X1 NAND2_1387 (.Y(N5604),.A(N3882),.B(N5112));
NAND2X1 NAND2_1388 (.Y(N5605),.A(N3879),.B(N5113));
NAND2X1 NAND2_1389 (.Y(N5631),.A(N5324),.B(N4653));
NAND2X1 NAND2_1390 (.Y(N5632),.A(N4463),.B(N5167));
NAND2X1 NAND2_1391 (.Y(N5640),.A(N4465),.B(N5168));
NAND2X1 NAND2_1392 (.Y(N5654),.A(N4467),.B(N5169));
NAND2X1 NAND2_1393 (.Y(N5670),.A(N4469),.B(N5170));
NAND2X1 NAND2_1394 (.Y(N5683),.A(N4471),.B(N5171));
NAND2X1 NAND2_1395 (.Y(N5690),.A(N4475),.B(N5172));
NAND2X1 NAND2_1396 (.Y(N5697),.A(N4477),.B(N5173));
NAND2X1 NAND2_1397 (.Y(N5707),.A(N4479),.B(N5174));
NAND2X1 NAND2_1398 (.Y(N5718),.A(N4481),.B(N5175));
NAND2X1 NAND2_1399 (.Y(N5728),.A(N4483),.B(N5176));
INVX1 NOT1_1400 (.Y(N5735),.A(N5177));
NAND2X1 NAND2_1401 (.Y(N5736),.A(N5179),.B(N4490));
NAND2X1 NAND2_1402 (.Y(N5740),.A(N5180),.B(N5181));
NAND2X1 NAND2_1403 (.Y(N5744),.A(N5182),.B(N5183));
NAND2X1 NAND2_1404 (.Y(N5747),.A(N5184),.B(N4496));
NAND2X1 NAND2_1405 (.Y(N5751),.A(N5185),.B(N5186));
NAND2X1 NAND2_1406 (.Y(N5755),.A(N5187),.B(N5188));
NAND2X1 NAND2_1407 (.Y(N5758),.A(N5189),.B(N4502));
NAND2X1 NAND2_1408 (.Y(N5762),.A(N5190),.B(N5191));
NAND2X1 NAND2_1409 (.Y(N5766),.A(N5192),.B(N5193));
INVX1 NOT1_1410 (.Y(N5769),.A(N4803));
INVX1 NOT1_1411 (.Y(N5770),.A(N4806));
NAND2X1 NAND2_1412 (.Y(N5771),.A(N4507),.B(N5196));
NAND2X1 NAND2_1413 (.Y(N5778),.A(N4509),.B(N5197));
NAND2X1 NAND2_1414 (.Y(N5789),.A(N4511),.B(N5198));
NAND2X1 NAND2_1415 (.Y(N5799),.A(N4513),.B(N5199));
NAND2X1 NAND2_1416 (.Y(N5807),.A(N4515),.B(N5200));
NAND2X1 NAND2_1417 (.Y(N5821),.A(N4517),.B(N5201));
NAND2X1 NAND2_1418 (.Y(N5837),.A(N4519),.B(N5202));
NAND2X1 NAND2_1419 (.Y(N5850),.A(N4521),.B(N5203));
NAND2X1 NAND2_1420 (.Y(N5856),.A(N4523),.B(N5204));
NAND2X1 NAND2_1421 (.Y(N5863),.A(N4525),.B(N5205));
NAND2X1 NAND2_1422 (.Y(N5870),.A(N4527),.B(N5206));
NAND2X1 NAND2_1423 (.Y(N5881),.A(N4529),.B(N5207));
NAND2X1 NAND2_1424 (.Y(N5892),.A(N4531),.B(N5208));
NAND2X1 NAND2_1425 (.Y(N5898),.A(N4533),.B(N5209));
NAND2X1 NAND2_1426 (.Y(N5905),.A(N4535),.B(N5210));
NAND2X1 NAND2_1427 (.Y(N5915),.A(N4537),.B(N5211));
NAND2X1 NAND2_1428 (.Y(N5926),.A(N4539),.B(N5212));
NAND2X1 NAND2_1429 (.Y(N5936),.A(N4541),.B(N5213));
INVX1 NOT1_1430 (.Y(N5943),.A(N4817));
NAND2X1 NAND2_1431 (.Y(N5944),.A(N4820),.B(N1931));
INVX1 NOT1_1432 (.Y(N5945),.A(N4820));
NAND2X1 NAND2_1433 (.Y(N5946),.A(N4823),.B(N1932));
INVX1 NOT1_1434 (.Y(N5947),.A(N4823));
NAND2X1 NAND2_1435 (.Y(N5948),.A(N4826),.B(N1933));
INVX1 NOT1_1436 (.Y(N5949),.A(N4826));
NAND2X1 NAND2_1437 (.Y(N5950),.A(N4829),.B(N1934));
INVX1 NOT1_1438 (.Y(N5951),.A(N4829));
NAND2X1 NAND2_1439 (.Y(N5952),.A(N4832),.B(N1935));
INVX1 NOT1_1440 (.Y(N5953),.A(N4832));
NAND2X1 NAND2_1441 (.Y(N5954),.A(N4835),.B(N1936));
INVX1 NOT1_1442 (.Y(N5955),.A(N4835));
NAND2X1 NAND2_1443 (.Y(N5956),.A(N4838),.B(N1937));
INVX1 NOT1_1444 (.Y(N5957),.A(N4838));
NAND2X1 NAND2_1445 (.Y(N5958),.A(N4841),.B(N1938));
INVX1 NOT1_1446 (.Y(N5959),.A(N4841));
AND2X1 AND2_1447 (.Y(N5960),.A(N2674),.B(N4769));
INVX1 NOT1_1448 (.Y(N5966),.A(N4844));
NAND2X1 NAND2_1449 (.Y(N5967),.A(N4847),.B(N1939));
INVX1 NOT1_1450 (.Y(N5968),.A(N4847));
NAND2X1 NAND2_1451 (.Y(N5969),.A(N4850),.B(N1940));
INVX1 NOT1_1452 (.Y(N5970),.A(N4850));
NAND2X1 NAND2_1453 (.Y(N5971),.A(N4853),.B(N1941));
INVX1 NOT1_1454 (.Y(N5972),.A(N4853));
NAND2X1 NAND2_1455 (.Y(N5973),.A(N4856),.B(N1942));
INVX1 NOT1_1456 (.Y(N5974),.A(N4856));
NAND2X1 NAND2_1457 (.Y(N5975),.A(N4859),.B(N1943));
INVX1 NOT1_1458 (.Y(N5976),.A(N4859));
NAND2X1 NAND2_1459 (.Y(N5977),.A(N4862),.B(N1944));
INVX1 NOT1_1460 (.Y(N5978),.A(N4862));
NAND2X1 NAND2_1461 (.Y(N5979),.A(N4865),.B(N1945));
INVX1 NOT1_1462 (.Y(N5980),.A(N4865));
AND2X1 AND2_1463 (.Y(N5981),.A(N2674),.B(N4769));
NAND2X1 NAND2_1464 (.Y(N5989),.A(N4868),.B(N1946));
INVX1 NOT1_1465 (.Y(N5990),.A(N4868));
NAND2X1 NAND2_1466 (.Y(N5991),.A(N5283),.B(N5284));
NAND2X1 NAND2_1467 (.Y(N5996),.A(N5285),.B(N5286));
NAND2X1 NAND2_1468 (.Y(N6000),.A(N5287),.B(N5288));
NAND2X1 NAND2_1469 (.Y(N6003),.A(N5289),.B(N5290));
NAND2X1 NAND2_1470 (.Y(N6009),.A(N5291),.B(N5292));
NAND2X1 NAND2_1471 (.Y(N6014),.A(N5293),.B(N5294));
NAND2X1 NAND2_1472 (.Y(N6018),.A(N5295),.B(N5296));
NAND2X1 NAND2_1473 (.Y(N6021),.A(N5297),.B(N5298));
NAND2X1 NAND2_1474 (.Y(N6022),.A(N5299),.B(N5300));
INVX1 NOT1_1475 (.Y(N6023),.A(N4874));
NAND2X1 NAND2_1476 (.Y(N6024),.A(N4874),.B(N4629));
INVX1 NOT1_1477 (.Y(N6025),.A(N4877));
NAND2X1 NAND2_1478 (.Y(N6026),.A(N4877),.B(N4631));
INVX1 NOT1_1479 (.Y(N6027),.A(N4880));
NAND2X1 NAND2_1480 (.Y(N6028),.A(N4880),.B(N4633));
INVX1 NOT1_1481 (.Y(N6029),.A(N4883));
NAND2X1 NAND2_1482 (.Y(N6030),.A(N4883),.B(N4636));
INVX1 NOT1_1483 (.Y(N6031),.A(N4886));
INVX1 NOT1_1484 (.Y(N6032),.A(N4889));
INVX1 NOT1_1485 (.Y(N6033),.A(N4892));
INVX1 NOT1_1486 (.Y(N6034),.A(N4895));
INVX1 NOT1_1487 (.Y(N6035),.A(N4898));
INVX1 NOT1_1488 (.Y(N6036),.A(N4901));
INVX1 NOT1_1489 (.Y(N6037),.A(N4904));
NAND2X1 NAND2_1490 (.Y(N6038),.A(N4904),.B(N4642));
INVX1 NOT1_1491 (.Y(N6039),.A(N4907));
INVX1 NOT1_1492 (.Y(N6040),.A(N4910));
NAND2X1 NAND2_1493 (.Y(N6041),.A(N5314),.B(N5315));
NAND2X1 NAND2_1494 (.Y(N6047),.A(N5316),.B(N5317));
NAND2X1 NAND2_1495 (.Y(N6052),.A(N5318),.B(N5319));
NAND2X1 NAND2_1496 (.Y(N6056),.A(N5320),.B(N5321));
NAND2X1 NAND2_1497 (.Y(N6059),.A(N5322),.B(N5323));
NAND2X1 NAND2_1498 (.Y(N6060),.A(N4913),.B(N1968));
INVX1 NOT1_1499 (.Y(N6061),.A(N4913));
NAND2X1 NAND2_1500 (.Y(N6062),.A(N4916),.B(N1969));
INVX1 NOT1_1501 (.Y(N6063),.A(N4916));
NAND2X1 NAND2_1502 (.Y(N6064),.A(N4919),.B(N1970));
INVX1 NOT1_1503 (.Y(N6065),.A(N4919));
NAND2X1 NAND2_1504 (.Y(N6066),.A(N4922),.B(N1971));
INVX1 NOT1_1505 (.Y(N6067),.A(N4922));
NAND2X1 NAND2_1506 (.Y(N6068),.A(N4925),.B(N1972));
INVX1 NOT1_1507 (.Y(N6069),.A(N4925));
NAND2X1 NAND2_1508 (.Y(N6070),.A(N4928),.B(N1973));
INVX1 NOT1_1509 (.Y(N6071),.A(N4928));
NAND2X1 NAND2_1510 (.Y(N6072),.A(N4931),.B(N1974));
INVX1 NOT1_1511 (.Y(N6073),.A(N4931));
NAND2X1 NAND2_1512 (.Y(N6074),.A(N4934),.B(N1975));
INVX1 NOT1_1513 (.Y(N6075),.A(N4934));
NAND2X1 NAND2_1514 (.Y(N6076),.A(N4937),.B(N1976));
INVX1 NOT1_1515 (.Y(N6077),.A(N4937));
INVX1 NOT1_1516 (.Y(N6078),.A(N4940));
NAND2X1 NAND2_1517 (.Y(N6079),.A(N5363),.B(N4694));
NAND2X1 NAND2_1518 (.Y(N6083),.A(N5364),.B(N5365));
NAND2X1 NAND2_1519 (.Y(N6087),.A(N5366),.B(N5367));
INVX1 NOT1_1520 (.Y(N6090),.A(N4943));
NAND2X1 NAND2_1521 (.Y(N6091),.A(N4943),.B(N4699));
INVX1 NOT1_1522 (.Y(N6092),.A(N4946));
INVX1 NOT1_1523 (.Y(N6093),.A(N4949));
INVX1 NOT1_1524 (.Y(N6094),.A(N4952));
INVX1 NOT1_1525 (.Y(N6095),.A(N4955));
INVX1 NOT1_1526 (.Y(N6096),.A(N4970));
NAND2X1 NAND2_1527 (.Y(N6097),.A(N4970),.B(N4700));
INVX1 NOT1_1528 (.Y(N6098),.A(N4973));
INVX1 NOT1_1529 (.Y(N6099),.A(N4976));
INVX1 NOT1_1530 (.Y(N6100),.A(N4979));
INVX1 NOT1_1531 (.Y(N6101),.A(N4982));
INVX1 NOT1_1532 (.Y(N6102),.A(N4997));
NAND2X1 NAND2_1533 (.Y(N6103),.A(N5000),.B(N2015));
INVX1 NOT1_1534 (.Y(N6104),.A(N5000));
NAND2X1 NAND2_1535 (.Y(N6105),.A(N5003),.B(N2016));
INVX1 NOT1_1536 (.Y(N6106),.A(N5003));
NAND2X1 NAND2_1537 (.Y(N6107),.A(N5006),.B(N2017));
INVX1 NOT1_1538 (.Y(N6108),.A(N5006));
NAND2X1 NAND2_1539 (.Y(N6109),.A(N5009),.B(N2018));
INVX1 NOT1_1540 (.Y(N6110),.A(N5009));
NAND2X1 NAND2_1541 (.Y(N6111),.A(N5012),.B(N2019));
INVX1 NOT1_1542 (.Y(N6112),.A(N5012));
NAND2X1 NAND2_1543 (.Y(N6113),.A(N5015),.B(N2020));
INVX1 NOT1_1544 (.Y(N6114),.A(N5015));
NAND2X1 NAND2_1545 (.Y(N6115),.A(N5018),.B(N2021));
INVX1 NOT1_1546 (.Y(N6116),.A(N5018));
NAND2X1 NAND2_1547 (.Y(N6117),.A(N5021),.B(N2022));
INVX1 NOT1_1548 (.Y(N6118),.A(N5021));
NAND2X1 NAND2_1549 (.Y(N6119),.A(N5024),.B(N2023));
INVX1 NOT1_1550 (.Y(N6120),.A(N5024));
INVX1 NOT1_1551 (.Y(N6121),.A(N5033));
NAND2X1 NAND2_1552 (.Y(N6122),.A(N5033),.B(N4743));
INVX1 NOT1_1553 (.Y(N6123),.A(N5036));
INVX1 NOT1_1554 (.Y(N6124),.A(N5039));
NAND2X1 NAND2_1555 (.Y(N6125),.A(N5042),.B(N4744));
INVX1 NOT1_1556 (.Y(N6126),.A(N5042));
NAND2X1 NAND2_1557 (.Y(N6127),.A(N5425),.B(N4746));
NAND2X1 NAND2_1558 (.Y(N6131),.A(N5426),.B(N5427));
INVX1 NOT1_1559 (.Y(N6135),.A(N5049));
NAND2X1 NAND2_1560 (.Y(N6136),.A(N5049),.B(N4749));
NAND2X1 NAND2_1561 (.Y(N6137),.A(N5429),.B(N4751));
NAND2X1 NAND2_1562 (.Y(N6141),.A(N5430),.B(N5431));
NAND2X1 NAND2_1563 (.Y(N6145),.A(N5432),.B(N5433));
INVX1 NOT1_1564 (.Y(N6148),.A(N5068));
INVX1 NOT1_1565 (.Y(N6149),.A(N5071));
INVX1 NOT1_1566 (.Y(N6150),.A(N5074));
INVX1 NOT1_1567 (.Y(N6151),.A(N5077));
INVX1 NOT1_1568 (.Y(N6152),.A(N5080));
INVX1 NOT1_1569 (.Y(N6153),.A(N5083));
INVX1 NOT1_1570 (.Y(N6154),.A(N5086));
INVX1 NOT1_1571 (.Y(N6155),.A(N5089));
INVX1 NOT1_1572 (.Y(N6156),.A(N5092));
NAND2X1 NAND2_1573 (.Y(N6157),.A(N5092),.B(N4761));
INVX1 NOT1_1574 (.Y(N6158),.A(N5095));
NAND2X1 NAND2_1575 (.Y(N6159),.A(N5095),.B(N4763));
INVX1 NOT1_1576 (.Y(N6160),.A(N5098));
NAND2X1 NAND2_1577 (.Y(N6161),.A(N5098),.B(N4765));
INVX1 NOT1_1578 (.Y(N6162),.A(N5101));
INVX1 NOT1_1579 (.Y(N6163),.A(N5104));
NAND2X1 NAND2_1580 (.Y(N6164),.A(N5107),.B(N4768));
INVX1 NOT1_1581 (.Y(N6165),.A(N5107));
NAND2X1 NAND2_1582 (.Y(N6166),.A(N5451),.B(N4776));
NAND2X1 NAND2_1583 (.Y(N6170),.A(N5452),.B(N5453));
NAND2X1 NAND2_1584 (.Y(N6174),.A(N5454),.B(N5455));
NAND2X1 NAND2_1585 (.Y(N6177),.A(N5456),.B(N5457));
INVX1 NOT1_1586 (.Y(N6181),.A(N5114));
INVX1 NOT1_1587 (.Y(N6182),.A(N5117));
INVX1 NOT1_1588 (.Y(N6183),.A(N5120));
INVX1 NOT1_1589 (.Y(N6184),.A(N5123));
INVX1 NOT1_1590 (.Y(N6185),.A(N5138));
NAND2X1 NAND2_1591 (.Y(N6186),.A(N5138),.B(N4783));
INVX1 NOT1_1592 (.Y(N6187),.A(N5141));
INVX1 NOT1_1593 (.Y(N6188),.A(N5144));
INVX1 NOT1_1594 (.Y(N6189),.A(N5147));
INVX1 NOT1_1595 (.Y(N6190),.A(N5150));
INVX1 NOT1_1596 (.Y(N6191),.A(N4784));
NAND2X1 NAND2_1597 (.Y(N6192),.A(N4784),.B(N2230));
INVX1 NOT1_1598 (.Y(N6193),.A(N4790));
NAND2X1 NAND2_1599 (.Y(N6194),.A(N4790),.B(N2765));
INVX1 NOT1_1600 (.Y(N6195),.A(N4796));
NAND2X1 NAND2_1601 (.Y(N6196),.A(N5476),.B(N5477));
NAND2X1 NAND2_1602 (.Y(N6199),.A(N5474),.B(N5475));
INVX1 NOT1_1603 (.Y(N6202),.A(N4810));
INVX1 NOT1_1604 (.Y(N6203),.A(N4814));
BUFX1 BUFF1_1605 (.Y(N6204),.A(N4769));
BUFX1 BUFF1_1606 (.Y(N6207),.A(N4555));
BUFX1 BUFF1_1607 (.Y(N6210),.A(N4769));
INVX1 NOT1_1608 (.Y(N6213),.A(N4871));
BUFX1 BUFF1_1609 (.Y(N6214),.A(N4586));
NOR2X1 NOR2_1610 (.Y(N6217),.A(N2674),.B(N4769));
BUFX1 BUFF1_1611 (.Y(N6220),.A(N4667));
INVX1 NOT1_1612 (.Y(N6223),.A(N4958));
INVX1 NOT1_1613 (.Y(N6224),.A(N4961));
INVX1 NOT1_1614 (.Y(N6225),.A(N4964));
INVX1 NOT1_1615 (.Y(N6226),.A(N4967));
INVX1 NOT1_1616 (.Y(N6227),.A(N4985));
INVX1 NOT1_1617 (.Y(N6228),.A(N4988));
INVX1 NOT1_1618 (.Y(N6229),.A(N4991));
INVX1 NOT1_1619 (.Y(N6230),.A(N4994));
INVX1 NOT1_1620 (.Y(N6231),.A(N5027));
BUFX1 BUFF1_1621 (.Y(N6232),.A(N4711));
INVX1 NOT1_1622 (.Y(N6235),.A(N5030));
BUFX1 BUFF1_1623 (.Y(N6236),.A(N4735));
INVX1 NOT1_1624 (.Y(N6239),.A(N5052));
INVX1 NOT1_1625 (.Y(N6240),.A(N5055));
INVX1 NOT1_1626 (.Y(N6241),.A(N5058));
INVX1 NOT1_1627 (.Y(N6242),.A(N5061));
NAND2X1 NAND2_1628 (.Y(N6243),.A(N5573),.B(N5574));
NAND2X1 NAND2_1629 (.Y(N6246),.A(N5571),.B(N5572));
NAND2X1 NAND2_1630 (.Y(N6249),.A(N5586),.B(N5587));
NAND2X1 NAND2_1631 (.Y(N6252),.A(N5584),.B(N5585));
INVX1 NOT1_1632 (.Y(N6255),.A(N5126));
INVX1 NOT1_1633 (.Y(N6256),.A(N5129));
INVX1 NOT1_1634 (.Y(N6257),.A(N5132));
INVX1 NOT1_1635 (.Y(N6258),.A(N5135));
INVX1 NOT1_1636 (.Y(N6259),.A(N5153));
INVX1 NOT1_1637 (.Y(N6260),.A(N5156));
INVX1 NOT1_1638 (.Y(N6261),.A(N5159));
INVX1 NOT1_1639 (.Y(N6262),.A(N5162));
NAND2X1 NAND2_1640 (.Y(N6263),.A(N5604),.B(N5605));
NAND2X1 NAND2_1641 (.Y(N6266),.A(N5602),.B(N5603));
NAND2X1 NAND2_1642 (.Y(N6540),.A(N1380),.B(N5945));
NAND2X1 NAND2_1643 (.Y(N6541),.A(N1383),.B(N5947));
NAND2X1 NAND2_1644 (.Y(N6542),.A(N1386),.B(N5949));
NAND2X1 NAND2_1645 (.Y(N6543),.A(N1389),.B(N5951));
NAND2X1 NAND2_1646 (.Y(N6544),.A(N1392),.B(N5953));
NAND2X1 NAND2_1647 (.Y(N6545),.A(N1395),.B(N5955));
NAND2X1 NAND2_1648 (.Y(N6546),.A(N1398),.B(N5957));
NAND2X1 NAND2_1649 (.Y(N6547),.A(N1401),.B(N5959));
NAND2X1 NAND2_1650 (.Y(N6555),.A(N1404),.B(N5968));
NAND2X1 NAND2_1651 (.Y(N6556),.A(N1407),.B(N5970));
NAND2X1 NAND2_1652 (.Y(N6557),.A(N1410),.B(N5972));
NAND2X1 NAND2_1653 (.Y(N6558),.A(N1413),.B(N5974));
NAND2X1 NAND2_1654 (.Y(N6559),.A(N1416),.B(N5976));
NAND2X1 NAND2_1655 (.Y(N6560),.A(N1419),.B(N5978));
NAND2X1 NAND2_1656 (.Y(N6561),.A(N1422),.B(N5980));
NAND2X1 NAND2_1657 (.Y(N6569),.A(N1425),.B(N5990));
NAND2X1 NAND2_1658 (.Y(N6594),.A(N3721),.B(N6023));
NAND2X1 NAND2_1659 (.Y(N6595),.A(N3724),.B(N6025));
NAND2X1 NAND2_1660 (.Y(N6596),.A(N3727),.B(N6027));
NAND2X1 NAND2_1661 (.Y(N6597),.A(N3730),.B(N6029));
NAND2X1 NAND2_1662 (.Y(N6598),.A(N4889),.B(N6031));
NAND2X1 NAND2_1663 (.Y(N6599),.A(N4886),.B(N6032));
NAND2X1 NAND2_1664 (.Y(N6600),.A(N4895),.B(N6033));
NAND2X1 NAND2_1665 (.Y(N6601),.A(N4892),.B(N6034));
NAND2X1 NAND2_1666 (.Y(N6602),.A(N4901),.B(N6035));
NAND2X1 NAND2_1667 (.Y(N6603),.A(N4898),.B(N6036));
NAND2X1 NAND2_1668 (.Y(N6604),.A(N3733),.B(N6037));
NAND2X1 NAND2_1669 (.Y(N6605),.A(N4910),.B(N6039));
NAND2X1 NAND2_1670 (.Y(N6606),.A(N4907),.B(N6040));
NAND2X1 NAND2_1671 (.Y(N6621),.A(N1434),.B(N6061));
NAND2X1 NAND2_1672 (.Y(N6622),.A(N1437),.B(N6063));
NAND2X1 NAND2_1673 (.Y(N6623),.A(N1440),.B(N6065));
NAND2X1 NAND2_1674 (.Y(N6624),.A(N1443),.B(N6067));
NAND2X1 NAND2_1675 (.Y(N6625),.A(N1446),.B(N6069));
NAND2X1 NAND2_1676 (.Y(N6626),.A(N1449),.B(N6071));
NAND2X1 NAND2_1677 (.Y(N6627),.A(N1452),.B(N6073));
NAND2X1 NAND2_1678 (.Y(N6628),.A(N1455),.B(N6075));
NAND2X1 NAND2_1679 (.Y(N6629),.A(N1458),.B(N6077));
NAND2X1 NAND2_1680 (.Y(N6639),.A(N3783),.B(N6090));
NAND2X1 NAND2_1681 (.Y(N6640),.A(N4949),.B(N6092));
NAND2X1 NAND2_1682 (.Y(N6641),.A(N4946),.B(N6093));
NAND2X1 NAND2_1683 (.Y(N6642),.A(N4955),.B(N6094));
NAND2X1 NAND2_1684 (.Y(N6643),.A(N4952),.B(N6095));
NAND2X1 NAND2_1685 (.Y(N6644),.A(N3786),.B(N6096));
NAND2X1 NAND2_1686 (.Y(N6645),.A(N4976),.B(N6098));
NAND2X1 NAND2_1687 (.Y(N6646),.A(N4973),.B(N6099));
NAND2X1 NAND2_1688 (.Y(N6647),.A(N4982),.B(N6100));
NAND2X1 NAND2_1689 (.Y(N6648),.A(N4979),.B(N6101));
NAND2X1 NAND2_1690 (.Y(N6649),.A(N1461),.B(N6104));
NAND2X1 NAND2_1691 (.Y(N6650),.A(N1464),.B(N6106));
NAND2X1 NAND2_1692 (.Y(N6651),.A(N1467),.B(N6108));
NAND2X1 NAND2_1693 (.Y(N6652),.A(N1470),.B(N6110));
NAND2X1 NAND2_1694 (.Y(N6653),.A(N1473),.B(N6112));
NAND2X1 NAND2_1695 (.Y(N6654),.A(N1476),.B(N6114));
NAND2X1 NAND2_1696 (.Y(N6655),.A(N1479),.B(N6116));
NAND2X1 NAND2_1697 (.Y(N6656),.A(N1482),.B(N6118));
NAND2X1 NAND2_1698 (.Y(N6657),.A(N1485),.B(N6120));
NAND2X1 NAND2_1699 (.Y(N6658),.A(N3789),.B(N6121));
NAND2X1 NAND2_1700 (.Y(N6659),.A(N5039),.B(N6123));
NAND2X1 NAND2_1701 (.Y(N6660),.A(N5036),.B(N6124));
NAND2X1 NAND2_1702 (.Y(N6661),.A(N3792),.B(N6126));
NAND2X1 NAND2_1703 (.Y(N6668),.A(N3816),.B(N6135));
NAND2X1 NAND2_1704 (.Y(N6677),.A(N5071),.B(N6148));
NAND2X1 NAND2_1705 (.Y(N6678),.A(N5068),.B(N6149));
NAND2X1 NAND2_1706 (.Y(N6679),.A(N5077),.B(N6150));
NAND2X1 NAND2_1707 (.Y(N6680),.A(N5074),.B(N6151));
NAND2X1 NAND2_1708 (.Y(N6681),.A(N5083),.B(N6152));
NAND2X1 NAND2_1709 (.Y(N6682),.A(N5080),.B(N6153));
NAND2X1 NAND2_1710 (.Y(N6683),.A(N5089),.B(N6154));
NAND2X1 NAND2_1711 (.Y(N6684),.A(N5086),.B(N6155));
NAND2X1 NAND2_1712 (.Y(N6685),.A(N3846),.B(N6156));
NAND2X1 NAND2_1713 (.Y(N6686),.A(N3849),.B(N6158));
NAND2X1 NAND2_1714 (.Y(N6687),.A(N3852),.B(N6160));
NAND2X1 NAND2_1715 (.Y(N6688),.A(N5104),.B(N6162));
NAND2X1 NAND2_1716 (.Y(N6689),.A(N5101),.B(N6163));
NAND2X1 NAND2_1717 (.Y(N6690),.A(N3855),.B(N6165));
NAND2X1 NAND2_1718 (.Y(N6702),.A(N5117),.B(N6181));
NAND2X1 NAND2_1719 (.Y(N6703),.A(N5114),.B(N6182));
NAND2X1 NAND2_1720 (.Y(N6704),.A(N5123),.B(N6183));
NAND2X1 NAND2_1721 (.Y(N6705),.A(N5120),.B(N6184));
NAND2X1 NAND2_1722 (.Y(N6706),.A(N3891),.B(N6185));
NAND2X1 NAND2_1723 (.Y(N6707),.A(N5144),.B(N6187));
NAND2X1 NAND2_1724 (.Y(N6708),.A(N5141),.B(N6188));
NAND2X1 NAND2_1725 (.Y(N6709),.A(N5150),.B(N6189));
NAND2X1 NAND2_1726 (.Y(N6710),.A(N5147),.B(N6190));
NAND2X1 NAND2_1727 (.Y(N6711),.A(N1708),.B(N6191));
NAND2X1 NAND2_1728 (.Y(N6712),.A(N2231),.B(N6193));
NAND2X1 NAND2_1729 (.Y(N6729),.A(N4961),.B(N6223));
NAND2X1 NAND2_1730 (.Y(N6730),.A(N4958),.B(N6224));
NAND2X1 NAND2_1731 (.Y(N6731),.A(N4967),.B(N6225));
NAND2X1 NAND2_1732 (.Y(N6732),.A(N4964),.B(N6226));
NAND2X1 NAND2_1733 (.Y(N6733),.A(N4988),.B(N6227));
NAND2X1 NAND2_1734 (.Y(N6734),.A(N4985),.B(N6228));
NAND2X1 NAND2_1735 (.Y(N6735),.A(N4994),.B(N6229));
NAND2X1 NAND2_1736 (.Y(N6736),.A(N4991),.B(N6230));
NAND2X1 NAND2_1737 (.Y(N6741),.A(N5055),.B(N6239));
NAND2X1 NAND2_1738 (.Y(N6742),.A(N5052),.B(N6240));
NAND2X1 NAND2_1739 (.Y(N6743),.A(N5061),.B(N6241));
NAND2X1 NAND2_1740 (.Y(N6744),.A(N5058),.B(N6242));
NAND2X1 NAND2_1741 (.Y(N6751),.A(N5129),.B(N6255));
NAND2X1 NAND2_1742 (.Y(N6752),.A(N5126),.B(N6256));
NAND2X1 NAND2_1743 (.Y(N6753),.A(N5135),.B(N6257));
NAND2X1 NAND2_1744 (.Y(N6754),.A(N5132),.B(N6258));
NAND2X1 NAND2_1745 (.Y(N6755),.A(N5156),.B(N6259));
NAND2X1 NAND2_1746 (.Y(N6756),.A(N5153),.B(N6260));
NAND2X1 NAND2_1747 (.Y(N6757),.A(N5162),.B(N6261));
NAND2X1 NAND2_1748 (.Y(N6758),.A(N5159),.B(N6262));
INVX1 NOT1_1749 (.Y(N6761),.A(N5892));
AND2X1 AND_tmp15 (.Y(ttmp15),.A(N5640),.B(N5632));
AND2X1 AND_tmp16 (.Y(ttmp16),.A(N5683),.B(ttmp15));
AND2X1 AND_tmp17 (.Y(ttmp17),.A(N5670),.B(ttmp16));
AND2X1 AND_tmp18 (.Y(N6762),.A(N5654),.B(ttmp17));
AND2X1 AND2_1751 (.Y(N6766),.A(N5632),.B(N3097));
AND2X1 AND_tmp19 (.Y(ttmp19),.A(N5632),.B(N3101));
AND2X1 AND_tmp20 (.Y(N6767),.A(N5640),.B(ttmp19));
AND2X1 AND_tmp21 (.Y(ttmp21),.A(N3107),.B(N5640));
AND2X1 AND_tmp22 (.Y(ttmp22),.A(N5654),.B(ttmp21));
AND2X1 AND_tmp23 (.Y(N6768),.A(N5632),.B(ttmp22));
AND2X1 AND_tmp24 (.Y(ttmp24),.A(N3114),.B(N5640));
AND2X1 AND_tmp25 (.Y(ttmp25),.A(N5670),.B(ttmp24));
AND2X1 AND_tmp26 (.Y(ttmp26),.A(N5654),.B(ttmp25));
AND2X1 AND_tmp27 (.Y(N6769),.A(N5632),.B(ttmp26));
AND2X1 AND2_1755 (.Y(N6770),.A(N5640),.B(N3101));
AND2X1 AND_tmp28 (.Y(ttmp28),.A(N3107),.B(N5640));
AND2X1 AND_tmp29 (.Y(N6771),.A(N5654),.B(ttmp28));
AND2X1 AND_tmp30 (.Y(ttmp30),.A(N3114),.B(N5640));
AND2X1 AND_tmp31 (.Y(ttmp31),.A(N5670),.B(ttmp30));
AND2X1 AND_tmp32 (.Y(N6772),.A(N5654),.B(ttmp31));
AND2X1 AND_tmp33 (.Y(ttmp33),.A(N5640),.B(N5670));
AND2X1 AND_tmp34 (.Y(ttmp34),.A(N5683),.B(ttmp33));
AND2X1 AND_tmp35 (.Y(N6773),.A(N5654),.B(ttmp34));
AND2X1 AND2_1759 (.Y(N6774),.A(N5640),.B(N3101));
AND2X1 AND_tmp36 (.Y(ttmp36),.A(N3107),.B(N5640));
AND2X1 AND_tmp37 (.Y(N6775),.A(N5654),.B(ttmp36));
AND2X1 AND_tmp38 (.Y(ttmp38),.A(N3114),.B(N5640));
AND2X1 AND_tmp39 (.Y(ttmp39),.A(N5670),.B(ttmp38));
AND2X1 AND_tmp40 (.Y(N6776),.A(N5654),.B(ttmp39));
AND2X1 AND2_1762 (.Y(N6777),.A(N5654),.B(N3107));
AND2X1 AND_tmp41 (.Y(ttmp41),.A(N5654),.B(N3114));
AND2X1 AND_tmp42 (.Y(N6778),.A(N5670),.B(ttmp41));
AND2X1 AND_tmp43 (.Y(ttmp43),.A(N5654),.B(N5670));
AND2X1 AND_tmp44 (.Y(N6779),.A(N5683),.B(ttmp43));
AND2X1 AND2_1765 (.Y(N6780),.A(N5654),.B(N3107));
AND2X1 AND_tmp45 (.Y(ttmp45),.A(N5654),.B(N3114));
AND2X1 AND_tmp46 (.Y(N6781),.A(N5670),.B(ttmp45));
AND2X1 AND2_1767 (.Y(N6782),.A(N5670),.B(N3114));
AND2X1 AND2_1768 (.Y(N6783),.A(N5683),.B(N5670));
AND2X1 AND_tmp47 (.Y(ttmp47),.A(N5690),.B(N5718));
AND2X1 AND_tmp48 (.Y(ttmp48),.A(N5697),.B(ttmp47));
AND2X1 AND_tmp49 (.Y(ttmp49),.A(N5728),.B(ttmp48));
AND2X1 AND_tmp50 (.Y(N6784),.A(N5707),.B(ttmp49));
AND2X1 AND2_1770 (.Y(N6787),.A(N5690),.B(N3137));
AND2X1 AND_tmp51 (.Y(ttmp51),.A(N5690),.B(N3140));
AND2X1 AND_tmp52 (.Y(N6788),.A(N5697),.B(ttmp51));
AND2X1 AND_tmp53 (.Y(ttmp53),.A(N3144),.B(N5697));
AND2X1 AND_tmp54 (.Y(ttmp54),.A(N5707),.B(ttmp53));
AND2X1 AND_tmp55 (.Y(N6789),.A(N5690),.B(ttmp54));
AND2X1 AND_tmp56 (.Y(ttmp56),.A(N3149),.B(N5697));
AND2X1 AND_tmp57 (.Y(ttmp57),.A(N5718),.B(ttmp56));
AND2X1 AND_tmp58 (.Y(ttmp58),.A(N5707),.B(ttmp57));
AND2X1 AND_tmp59 (.Y(N6790),.A(N5690),.B(ttmp58));
AND2X1 AND2_1774 (.Y(N6791),.A(N5697),.B(N3140));
AND2X1 AND_tmp60 (.Y(ttmp60),.A(N3144),.B(N5697));
AND2X1 AND_tmp61 (.Y(N6792),.A(N5707),.B(ttmp60));
AND2X1 AND_tmp62 (.Y(ttmp62),.A(N3149),.B(N5697));
AND2X1 AND_tmp63 (.Y(ttmp63),.A(N5718),.B(ttmp62));
AND2X1 AND_tmp64 (.Y(N6793),.A(N5707),.B(ttmp63));
AND2X1 AND2_1777 (.Y(N6794),.A(N3144),.B(N5707));
AND2X1 AND_tmp65 (.Y(ttmp65),.A(N5707),.B(N3149));
AND2X1 AND_tmp66 (.Y(N6795),.A(N5718),.B(ttmp65));
AND2X1 AND2_1779 (.Y(N6796),.A(N5718),.B(N3149));
INVX1 NOT1_1780 (.Y(N6797),.A(N5736));
INVX1 NOT1_1781 (.Y(N6800),.A(N5740));
INVX1 NOT1_1782 (.Y(N6803),.A(N5747));
INVX1 NOT1_1783 (.Y(N6806),.A(N5751));
INVX1 NOT1_1784 (.Y(N6809),.A(N5758));
INVX1 NOT1_1785 (.Y(N6812),.A(N5762));
BUFX1 BUFF1_1786 (.Y(N6815),.A(N5744));
BUFX1 BUFF1_1787 (.Y(N6818),.A(N5744));
BUFX1 BUFF1_1788 (.Y(N6821),.A(N5755));
BUFX1 BUFF1_1789 (.Y(N6824),.A(N5755));
BUFX1 BUFF1_1790 (.Y(N6827),.A(N5766));
BUFX1 BUFF1_1791 (.Y(N6830),.A(N5766));
AND2X1 AND_tmp67 (.Y(ttmp67),.A(N5778),.B(N5771));
AND2X1 AND_tmp68 (.Y(ttmp68),.A(N5850),.B(ttmp67));
AND2X1 AND_tmp69 (.Y(N6833),.A(N5789),.B(ttmp68));
AND2X1 AND2_1793 (.Y(N6836),.A(N5771),.B(N3169));
AND2X1 AND_tmp70 (.Y(ttmp70),.A(N5771),.B(N3173));
AND2X1 AND_tmp71 (.Y(N6837),.A(N5778),.B(ttmp70));
AND2X1 AND_tmp72 (.Y(ttmp72),.A(N3178),.B(N5778));
AND2X1 AND_tmp73 (.Y(ttmp73),.A(N5789),.B(ttmp72));
AND2X1 AND_tmp74 (.Y(N6838),.A(N5771),.B(ttmp73));
AND2X1 AND2_1796 (.Y(N6839),.A(N5778),.B(N3173));
AND2X1 AND_tmp75 (.Y(ttmp75),.A(N3178),.B(N5778));
AND2X1 AND_tmp76 (.Y(N6840),.A(N5789),.B(ttmp75));
AND2X1 AND_tmp77 (.Y(ttmp77),.A(N5789),.B(N5778));
AND2X1 AND_tmp78 (.Y(N6841),.A(N5850),.B(ttmp77));
AND2X1 AND2_1799 (.Y(N6842),.A(N5778),.B(N3173));
AND2X1 AND_tmp79 (.Y(ttmp79),.A(N3178),.B(N5778));
AND2X1 AND_tmp80 (.Y(N6843),.A(N5789),.B(ttmp79));
AND2X1 AND2_1801 (.Y(N6844),.A(N5789),.B(N3178));
AND2X1 AND_tmp81 (.Y(ttmp81),.A(N5807),.B(N5799));
AND2X1 AND_tmp82 (.Y(ttmp82),.A(N5856),.B(ttmp81));
AND2X1 AND_tmp83 (.Y(ttmp83),.A(N5837),.B(ttmp82));
AND2X1 AND_tmp84 (.Y(N6845),.A(N5821),.B(ttmp83));
AND2X1 AND2_1803 (.Y(N6848),.A(N5799),.B(N3185));
AND2X1 AND_tmp85 (.Y(ttmp85),.A(N5799),.B(N3189));
AND2X1 AND_tmp86 (.Y(N6849),.A(N5807),.B(ttmp85));
AND2X1 AND_tmp87 (.Y(ttmp87),.A(N3195),.B(N5807));
AND2X1 AND_tmp88 (.Y(ttmp88),.A(N5821),.B(ttmp87));
AND2X1 AND_tmp89 (.Y(N6850),.A(N5799),.B(ttmp88));
AND2X1 AND_tmp90 (.Y(ttmp90),.A(N3202),.B(N5807));
AND2X1 AND_tmp91 (.Y(ttmp91),.A(N5837),.B(ttmp90));
AND2X1 AND_tmp92 (.Y(ttmp92),.A(N5821),.B(ttmp91));
AND2X1 AND_tmp93 (.Y(N6851),.A(N5799),.B(ttmp92));
AND2X1 AND2_1807 (.Y(N6852),.A(N5807),.B(N3189));
AND2X1 AND_tmp94 (.Y(ttmp94),.A(N3195),.B(N5807));
AND2X1 AND_tmp95 (.Y(N6853),.A(N5821),.B(ttmp94));
AND2X1 AND_tmp96 (.Y(ttmp96),.A(N3202),.B(N5807));
AND2X1 AND_tmp97 (.Y(ttmp97),.A(N5837),.B(ttmp96));
AND2X1 AND_tmp98 (.Y(N6854),.A(N5821),.B(ttmp97));
AND2X1 AND_tmp99 (.Y(ttmp99),.A(N5807),.B(N5837));
AND2X1 AND_tmp100 (.Y(ttmp100),.A(N5856),.B(ttmp99));
AND2X1 AND_tmp101 (.Y(N6855),.A(N5821),.B(ttmp100));
AND2X1 AND2_1811 (.Y(N6856),.A(N5807),.B(N3189));
AND2X1 AND_tmp102 (.Y(ttmp102),.A(N3195),.B(N5807));
AND2X1 AND_tmp103 (.Y(N6857),.A(N5821),.B(ttmp102));
AND2X1 AND_tmp104 (.Y(ttmp104),.A(N3202),.B(N5807));
AND2X1 AND_tmp105 (.Y(ttmp105),.A(N5837),.B(ttmp104));
AND2X1 AND_tmp106 (.Y(N6858),.A(N5821),.B(ttmp105));
AND2X1 AND2_1814 (.Y(N6859),.A(N5821),.B(N3195));
AND2X1 AND_tmp107 (.Y(ttmp107),.A(N5821),.B(N3202));
AND2X1 AND_tmp108 (.Y(N6860),.A(N5837),.B(ttmp107));
AND2X1 AND_tmp109 (.Y(ttmp109),.A(N5821),.B(N5837));
AND2X1 AND_tmp110 (.Y(N6861),.A(N5856),.B(ttmp109));
AND2X1 AND2_1817 (.Y(N6862),.A(N5821),.B(N3195));
AND2X1 AND_tmp111 (.Y(ttmp111),.A(N5821),.B(N3202));
AND2X1 AND_tmp112 (.Y(N6863),.A(N5837),.B(ttmp111));
AND2X1 AND2_1819 (.Y(N6864),.A(N5837),.B(N3202));
AND2X1 AND2_1820 (.Y(N6865),.A(N5850),.B(N5789));
AND2X1 AND2_1821 (.Y(N6866),.A(N5856),.B(N5837));
AND2X1 AND_tmp113 (.Y(ttmp113),.A(N5881),.B(N5863));
AND2X1 AND_tmp114 (.Y(ttmp114),.A(N5870),.B(ttmp113));
AND2X1 AND_tmp115 (.Y(N6867),.A(N5892),.B(ttmp114));
AND2X1 AND2_1823 (.Y(N6870),.A(N5863),.B(N3211));
AND2X1 AND_tmp116 (.Y(ttmp116),.A(N5863),.B(N3215));
AND2X1 AND_tmp117 (.Y(N6871),.A(N5870),.B(ttmp116));
AND2X1 AND_tmp118 (.Y(ttmp118),.A(N3221),.B(N5870));
AND2X1 AND_tmp119 (.Y(ttmp119),.A(N5881),.B(ttmp118));
AND2X1 AND_tmp120 (.Y(N6872),.A(N5863),.B(ttmp119));
AND2X1 AND2_1826 (.Y(N6873),.A(N5870),.B(N3215));
AND2X1 AND_tmp121 (.Y(ttmp121),.A(N3221),.B(N5870));
AND2X1 AND_tmp122 (.Y(N6874),.A(N5881),.B(ttmp121));
AND2X1 AND_tmp123 (.Y(ttmp123),.A(N5881),.B(N5870));
AND2X1 AND_tmp124 (.Y(N6875),.A(N5892),.B(ttmp123));
AND2X1 AND2_1829 (.Y(N6876),.A(N5870),.B(N3215));
AND2X1 AND_tmp125 (.Y(ttmp125),.A(N5881),.B(N5870));
AND2X1 AND_tmp126 (.Y(N6877),.A(N3221),.B(ttmp125));
AND2X1 AND2_1831 (.Y(N6878),.A(N5881),.B(N3221));
AND2X1 AND2_1832 (.Y(N6879),.A(N5892),.B(N5881));
AND2X1 AND2_1833 (.Y(N6880),.A(N5881),.B(N3221));
AND2X1 AND_tmp127 (.Y(ttmp127),.A(N5898),.B(N5926));
AND2X1 AND_tmp128 (.Y(ttmp128),.A(N5905),.B(ttmp127));
AND2X1 AND_tmp129 (.Y(ttmp129),.A(N5936),.B(ttmp128));
AND2X1 AND_tmp130 (.Y(N6881),.A(N5915),.B(ttmp129));
AND2X1 AND2_1835 (.Y(N6884),.A(N5898),.B(N3229));
AND2X1 AND_tmp131 (.Y(ttmp131),.A(N5898),.B(N3232));
AND2X1 AND_tmp132 (.Y(N6885),.A(N5905),.B(ttmp131));
AND2X1 AND_tmp133 (.Y(ttmp133),.A(N3236),.B(N5905));
AND2X1 AND_tmp134 (.Y(ttmp134),.A(N5915),.B(ttmp133));
AND2X1 AND_tmp135 (.Y(N6886),.A(N5898),.B(ttmp134));
AND2X1 AND_tmp136 (.Y(ttmp136),.A(N3241),.B(N5905));
AND2X1 AND_tmp137 (.Y(ttmp137),.A(N5926),.B(ttmp136));
AND2X1 AND_tmp138 (.Y(ttmp138),.A(N5915),.B(ttmp137));
AND2X1 AND_tmp139 (.Y(N6887),.A(N5898),.B(ttmp138));
AND2X1 AND2_1839 (.Y(N6888),.A(N5905),.B(N3232));
AND2X1 AND_tmp140 (.Y(ttmp140),.A(N3236),.B(N5905));
AND2X1 AND_tmp141 (.Y(N6889),.A(N5915),.B(ttmp140));
AND2X1 AND_tmp142 (.Y(ttmp142),.A(N3241),.B(N5905));
AND2X1 AND_tmp143 (.Y(ttmp143),.A(N5926),.B(ttmp142));
AND2X1 AND_tmp144 (.Y(N6890),.A(N5915),.B(ttmp143));
AND2X1 AND2_1842 (.Y(N6891),.A(N3236),.B(N5915));
AND2X1 AND_tmp145 (.Y(ttmp145),.A(N5915),.B(N3241));
AND2X1 AND_tmp146 (.Y(N6892),.A(N5926),.B(ttmp145));
AND2X1 AND2_1844 (.Y(N6893),.A(N5926),.B(N3241));
NAND2X1 NAND2_1845 (.Y(N6894),.A(N5944),.B(N6540));
NAND2X1 NAND2_1846 (.Y(N6901),.A(N5946),.B(N6541));
NAND2X1 NAND2_1847 (.Y(N6912),.A(N5948),.B(N6542));
NAND2X1 NAND2_1848 (.Y(N6923),.A(N5950),.B(N6543));
NAND2X1 NAND2_1849 (.Y(N6929),.A(N5952),.B(N6544));
NAND2X1 NAND2_1850 (.Y(N6936),.A(N5954),.B(N6545));
NAND2X1 NAND2_1851 (.Y(N6946),.A(N5956),.B(N6546));
NAND2X1 NAND2_1852 (.Y(N6957),.A(N5958),.B(N6547));
NAND2X1 NAND2_1853 (.Y(N6967),.A(N6204),.B(N4575));
INVX1 NOT1_1854 (.Y(N6968),.A(N6204));
INVX1 NOT1_1855 (.Y(N6969),.A(N6207));
NAND2X1 NAND2_1856 (.Y(N6970),.A(N5967),.B(N6555));
NAND2X1 NAND2_1857 (.Y(N6977),.A(N5969),.B(N6556));
NAND2X1 NAND2_1858 (.Y(N6988),.A(N5971),.B(N6557));
NAND2X1 NAND2_1859 (.Y(N6998),.A(N5973),.B(N6558));
NAND2X1 NAND2_1860 (.Y(N7006),.A(N5975),.B(N6559));
NAND2X1 NAND2_1861 (.Y(N7020),.A(N5977),.B(N6560));
NAND2X1 NAND2_1862 (.Y(N7036),.A(N5979),.B(N6561));
NAND2X1 NAND2_1863 (.Y(N7049),.A(N5989),.B(N6569));
NAND2X1 NAND2_1864 (.Y(N7055),.A(N6210),.B(N4610));
INVX1 NOT1_1865 (.Y(N7056),.A(N6210));
AND2X1 AND_tmp147 (.Y(ttmp147),.A(N5996),.B(N5991));
AND2X1 AND_tmp148 (.Y(ttmp148),.A(N6021),.B(ttmp147));
AND2X1 AND_tmp149 (.Y(N7057),.A(N6000),.B(ttmp148));
AND2X1 AND2_1867 (.Y(N7060),.A(N5991),.B(N3362));
AND2X1 AND_tmp150 (.Y(ttmp150),.A(N5991),.B(N3363));
AND2X1 AND_tmp151 (.Y(N7061),.A(N5996),.B(ttmp150));
AND2X1 AND_tmp152 (.Y(ttmp152),.A(N3364),.B(N5996));
AND2X1 AND_tmp153 (.Y(ttmp153),.A(N6000),.B(ttmp152));
AND2X1 AND_tmp154 (.Y(N7062),.A(N5991),.B(ttmp153));
AND2X1 AND_tmp155 (.Y(ttmp155),.A(N6009),.B(N6003));
AND2X1 AND_tmp156 (.Y(ttmp156),.A(N6022),.B(ttmp155));
AND2X1 AND_tmp157 (.Y(ttmp157),.A(N6018),.B(ttmp156));
AND2X1 AND_tmp158 (.Y(N7063),.A(N6014),.B(ttmp157));
AND2X1 AND2_1871 (.Y(N7064),.A(N6003),.B(N3366));
AND2X1 AND_tmp159 (.Y(ttmp159),.A(N6003),.B(N3367));
AND2X1 AND_tmp160 (.Y(N7065),.A(N6009),.B(ttmp159));
AND2X1 AND_tmp161 (.Y(ttmp161),.A(N3368),.B(N6009));
AND2X1 AND_tmp162 (.Y(ttmp162),.A(N6014),.B(ttmp161));
AND2X1 AND_tmp163 (.Y(N7066),.A(N6003),.B(ttmp162));
AND2X1 AND_tmp164 (.Y(ttmp164),.A(N3369),.B(N6009));
AND2X1 AND_tmp165 (.Y(ttmp165),.A(N6018),.B(ttmp164));
AND2X1 AND_tmp166 (.Y(ttmp166),.A(N6014),.B(ttmp165));
AND2X1 AND_tmp167 (.Y(N7067),.A(N6003),.B(ttmp166));
NAND2X1 NAND2_1875 (.Y(N7068),.A(N6594),.B(N6024));
NAND2X1 NAND2_1876 (.Y(N7073),.A(N6595),.B(N6026));
NAND2X1 NAND2_1877 (.Y(N7077),.A(N6596),.B(N6028));
NAND2X1 NAND2_1878 (.Y(N7080),.A(N6597),.B(N6030));
NAND2X1 NAND2_1879 (.Y(N7086),.A(N6598),.B(N6599));
NAND2X1 NAND2_1880 (.Y(N7091),.A(N6600),.B(N6601));
NAND2X1 NAND2_1881 (.Y(N7095),.A(N6602),.B(N6603));
NAND2X1 NAND2_1882 (.Y(N7098),.A(N6604),.B(N6038));
NAND2X1 NAND2_1883 (.Y(N7099),.A(N6605),.B(N6606));
AND2X1 AND_tmp168 (.Y(ttmp168),.A(N6047),.B(N6041));
AND2X1 AND_tmp169 (.Y(ttmp169),.A(N6059),.B(ttmp168));
AND2X1 AND_tmp170 (.Y(ttmp170),.A(N6056),.B(ttmp169));
AND2X1 AND_tmp171 (.Y(N7100),.A(N6052),.B(ttmp170));
AND2X1 AND2_1885 (.Y(N7103),.A(N6041),.B(N3371));
AND2X1 AND_tmp172 (.Y(ttmp172),.A(N6041),.B(N3372));
AND2X1 AND_tmp173 (.Y(N7104),.A(N6047),.B(ttmp172));
AND2X1 AND_tmp174 (.Y(ttmp174),.A(N3373),.B(N6047));
AND2X1 AND_tmp175 (.Y(ttmp175),.A(N6052),.B(ttmp174));
AND2X1 AND_tmp176 (.Y(N7105),.A(N6041),.B(ttmp175));
AND2X1 AND_tmp177 (.Y(ttmp177),.A(N3374),.B(N6047));
AND2X1 AND_tmp178 (.Y(ttmp178),.A(N6056),.B(ttmp177));
AND2X1 AND_tmp179 (.Y(ttmp179),.A(N6052),.B(ttmp178));
AND2X1 AND_tmp180 (.Y(N7106),.A(N6041),.B(ttmp179));
NAND2X1 NAND2_1889 (.Y(N7107),.A(N6060),.B(N6621));
NAND2X1 NAND2_1890 (.Y(N7114),.A(N6062),.B(N6622));
NAND2X1 NAND2_1891 (.Y(N7125),.A(N6064),.B(N6623));
NAND2X1 NAND2_1892 (.Y(N7136),.A(N6066),.B(N6624));
NAND2X1 NAND2_1893 (.Y(N7142),.A(N6068),.B(N6625));
NAND2X1 NAND2_1894 (.Y(N7149),.A(N6070),.B(N6626));
NAND2X1 NAND2_1895 (.Y(N7159),.A(N6072),.B(N6627));
NAND2X1 NAND2_1896 (.Y(N7170),.A(N6074),.B(N6628));
NAND2X1 NAND2_1897 (.Y(N7180),.A(N6076),.B(N6629));
INVX1 NOT1_1898 (.Y(N7187),.A(N6220));
INVX1 NOT1_1899 (.Y(N7188),.A(N6079));
INVX1 NOT1_1900 (.Y(N7191),.A(N6083));
NAND2X1 NAND2_1901 (.Y(N7194),.A(N6639),.B(N6091));
NAND2X1 NAND2_1902 (.Y(N7198),.A(N6640),.B(N6641));
NAND2X1 NAND2_1903 (.Y(N7202),.A(N6642),.B(N6643));
NAND2X1 NAND2_1904 (.Y(N7205),.A(N6644),.B(N6097));
NAND2X1 NAND2_1905 (.Y(N7209),.A(N6645),.B(N6646));
NAND2X1 NAND2_1906 (.Y(N7213),.A(N6647),.B(N6648));
BUFX1 BUFF1_1907 (.Y(N7216),.A(N6087));
BUFX1 BUFF1_1908 (.Y(N7219),.A(N6087));
NAND2X1 NAND2_1909 (.Y(N7222),.A(N6103),.B(N6649));
NAND2X1 NAND2_1910 (.Y(N7229),.A(N6105),.B(N6650));
NAND2X1 NAND2_1911 (.Y(N7240),.A(N6107),.B(N6651));
NAND2X1 NAND2_1912 (.Y(N7250),.A(N6109),.B(N6652));
NAND2X1 NAND2_1913 (.Y(N7258),.A(N6111),.B(N6653));
NAND2X1 NAND2_1914 (.Y(N7272),.A(N6113),.B(N6654));
NAND2X1 NAND2_1915 (.Y(N7288),.A(N6115),.B(N6655));
NAND2X1 NAND2_1916 (.Y(N7301),.A(N6117),.B(N6656));
NAND2X1 NAND2_1917 (.Y(N7307),.A(N6119),.B(N6657));
NAND2X1 NAND2_1918 (.Y(N7314),.A(N6658),.B(N6122));
NAND2X1 NAND2_1919 (.Y(N7318),.A(N6659),.B(N6660));
NAND2X1 NAND2_1920 (.Y(N7322),.A(N6125),.B(N6661));
INVX1 NOT1_1921 (.Y(N7325),.A(N6127));
INVX1 NOT1_1922 (.Y(N7328),.A(N6131));
NAND2X1 NAND2_1923 (.Y(N7331),.A(N6668),.B(N6136));
INVX1 NOT1_1924 (.Y(N7334),.A(N6137));
INVX1 NOT1_1925 (.Y(N7337),.A(N6141));
BUFX1 BUFF1_1926 (.Y(N7340),.A(N6145));
BUFX1 BUFF1_1927 (.Y(N7343),.A(N6145));
NAND2X1 NAND2_1928 (.Y(N7346),.A(N6677),.B(N6678));
NAND2X1 NAND2_1929 (.Y(N7351),.A(N6679),.B(N6680));
NAND2X1 NAND2_1930 (.Y(N7355),.A(N6681),.B(N6682));
NAND2X1 NAND2_1931 (.Y(N7358),.A(N6683),.B(N6684));
NAND2X1 NAND2_1932 (.Y(N7364),.A(N6685),.B(N6157));
NAND2X1 NAND2_1933 (.Y(N7369),.A(N6686),.B(N6159));
NAND2X1 NAND2_1934 (.Y(N7373),.A(N6687),.B(N6161));
NAND2X1 NAND2_1935 (.Y(N7376),.A(N6688),.B(N6689));
NAND2X1 NAND2_1936 (.Y(N7377),.A(N6164),.B(N6690));
INVX1 NOT1_1937 (.Y(N7378),.A(N6166));
INVX1 NOT1_1938 (.Y(N7381),.A(N6170));
INVX1 NOT1_1939 (.Y(N7384),.A(N6177));
NAND2X1 NAND2_1940 (.Y(N7387),.A(N6702),.B(N6703));
NAND2X1 NAND2_1941 (.Y(N7391),.A(N6704),.B(N6705));
NAND2X1 NAND2_1942 (.Y(N7394),.A(N6706),.B(N6186));
NAND2X1 NAND2_1943 (.Y(N7398),.A(N6707),.B(N6708));
NAND2X1 NAND2_1944 (.Y(N7402),.A(N6709),.B(N6710));
BUFX1 BUFF1_1945 (.Y(N7405),.A(N6174));
BUFX1 BUFF1_1946 (.Y(N7408),.A(N6174));
BUFX1 BUFF1_1947 (.Y(N7411),.A(N5936));
BUFX1 BUFF1_1948 (.Y(N7414),.A(N5898));
BUFX1 BUFF1_1949 (.Y(N7417),.A(N5905));
BUFX1 BUFF1_1950 (.Y(N7420),.A(N5915));
BUFX1 BUFF1_1951 (.Y(N7423),.A(N5926));
BUFX1 BUFF1_1952 (.Y(N7426),.A(N5728));
BUFX1 BUFF1_1953 (.Y(N7429),.A(N5690));
BUFX1 BUFF1_1954 (.Y(N7432),.A(N5697));
BUFX1 BUFF1_1955 (.Y(N7435),.A(N5707));
BUFX1 BUFF1_1956 (.Y(N7438),.A(N5718));
NAND2X1 NAND2_1957 (.Y(N7441),.A(N6192),.B(N6711));
NAND2X1 NAND2_1958 (.Y(N7444),.A(N6194),.B(N6712));
BUFX1 BUFF1_1959 (.Y(N7447),.A(N5683));
BUFX1 BUFF1_1960 (.Y(N7450),.A(N5670));
BUFX1 BUFF1_1961 (.Y(N7453),.A(N5632));
BUFX1 BUFF1_1962 (.Y(N7456),.A(N5654));
BUFX1 BUFF1_1963 (.Y(N7459),.A(N5640));
BUFX1 BUFF1_1964 (.Y(N7462),.A(N5640));
BUFX1 BUFF1_1965 (.Y(N7465),.A(N5683));
BUFX1 BUFF1_1966 (.Y(N7468),.A(N5670));
BUFX1 BUFF1_1967 (.Y(N7471),.A(N5632));
BUFX1 BUFF1_1968 (.Y(N7474),.A(N5654));
INVX1 NOT1_1969 (.Y(N7477),.A(N6196));
INVX1 NOT1_1970 (.Y(N7478),.A(N6199));
BUFX1 BUFF1_1971 (.Y(N7479),.A(N5850));
BUFX1 BUFF1_1972 (.Y(N7482),.A(N5789));
BUFX1 BUFF1_1973 (.Y(N7485),.A(N5771));
BUFX1 BUFF1_1974 (.Y(N7488),.A(N5778));
BUFX1 BUFF1_1975 (.Y(N7491),.A(N5850));
BUFX1 BUFF1_1976 (.Y(N7494),.A(N5789));
BUFX1 BUFF1_1977 (.Y(N7497),.A(N5771));
BUFX1 BUFF1_1978 (.Y(N7500),.A(N5778));
BUFX1 BUFF1_1979 (.Y(N7503),.A(N5856));
BUFX1 BUFF1_1980 (.Y(N7506),.A(N5837));
BUFX1 BUFF1_1981 (.Y(N7509),.A(N5799));
BUFX1 BUFF1_1982 (.Y(N7512),.A(N5821));
BUFX1 BUFF1_1983 (.Y(N7515),.A(N5807));
BUFX1 BUFF1_1984 (.Y(N7518),.A(N5807));
BUFX1 BUFF1_1985 (.Y(N7521),.A(N5856));
BUFX1 BUFF1_1986 (.Y(N7524),.A(N5837));
BUFX1 BUFF1_1987 (.Y(N7527),.A(N5799));
BUFX1 BUFF1_1988 (.Y(N7530),.A(N5821));
BUFX1 BUFF1_1989 (.Y(N7533),.A(N5863));
BUFX1 BUFF1_1990 (.Y(N7536),.A(N5863));
BUFX1 BUFF1_1991 (.Y(N7539),.A(N5870));
BUFX1 BUFF1_1992 (.Y(N7542),.A(N5870));
BUFX1 BUFF1_1993 (.Y(N7545),.A(N5881));
BUFX1 BUFF1_1994 (.Y(N7548),.A(N5881));
INVX1 NOT1_1995 (.Y(N7551),.A(N6214));
INVX1 NOT1_1996 (.Y(N7552),.A(N6217));
BUFX1 BUFF1_1997 (.Y(N7553),.A(N5981));
INVX1 NOT1_1998 (.Y(N7556),.A(N6249));
INVX1 NOT1_1999 (.Y(N7557),.A(N6252));
INVX1 NOT1_2000 (.Y(N7558),.A(N6243));
INVX1 NOT1_2001 (.Y(N7559),.A(N6246));
NAND2X1 NAND2_2002 (.Y(N7560),.A(N6731),.B(N6732));
NAND2X1 NAND2_2003 (.Y(N7563),.A(N6729),.B(N6730));
NAND2X1 NAND2_2004 (.Y(N7566),.A(N6735),.B(N6736));
NAND2X1 NAND2_2005 (.Y(N7569),.A(N6733),.B(N6734));
INVX1 NOT1_2006 (.Y(N7572),.A(N6232));
INVX1 NOT1_2007 (.Y(N7573),.A(N6236));
NAND2X1 NAND2_2008 (.Y(N7574),.A(N6743),.B(N6744));
NAND2X1 NAND2_2009 (.Y(N7577),.A(N6741),.B(N6742));
INVX1 NOT1_2010 (.Y(N7580),.A(N6263));
INVX1 NOT1_2011 (.Y(N7581),.A(N6266));
NAND2X1 NAND2_2012 (.Y(N7582),.A(N6753),.B(N6754));
NAND2X1 NAND2_2013 (.Y(N7585),.A(N6751),.B(N6752));
NAND2X1 NAND2_2014 (.Y(N7588),.A(N6757),.B(N6758));
NAND2X1 NAND2_2015 (.Y(N7591),.A(N6755),.B(N6756));
OR2X1 OR_tmp181 (.Y(ttmp181),.A(N6768),.B(N6769));
OR2X1 OR_tmp182 (.Y(ttmp182),.A(N3096),.B(ttmp181));
OR2X1 OR_tmp183 (.Y(ttmp183),.A(N6766),.B(ttmp182));
OR2X1 OR_tmp184 (.Y(N7609),.A(N6767),.B(ttmp183));
OR2X1 OR2_2017 (.Y(N7613),.A(N3107),.B(N6782));
OR2X1 OR_tmp185 (.Y(ttmp185),.A(N6789),.B(N6790));
OR2X1 OR_tmp186 (.Y(ttmp186),.A(N3136),.B(ttmp185));
OR2X1 OR_tmp187 (.Y(ttmp187),.A(N6787),.B(ttmp186));
OR2X1 OR_tmp188 (.Y(N7620),.A(N6788),.B(ttmp187));
OR2X1 OR_tmp189 (.Y(ttmp189),.A(N6837),.B(N6838));
OR2X1 OR_tmp190 (.Y(ttmp190),.A(N3168),.B(ttmp189));
OR2X1 OR_tmp191 (.Y(N7649),.A(N6836),.B(ttmp190));
OR2X1 OR2_2020 (.Y(N7650),.A(N3173),.B(N6844));
OR2X1 OR_tmp192 (.Y(ttmp192),.A(N6850),.B(N6851));
OR2X1 OR_tmp193 (.Y(ttmp193),.A(N3184),.B(ttmp192));
OR2X1 OR_tmp194 (.Y(ttmp194),.A(N6848),.B(ttmp193));
OR2X1 OR_tmp195 (.Y(N7655),.A(N6849),.B(ttmp194));
OR2X1 OR2_2022 (.Y(N7659),.A(N3195),.B(N6864));
OR2X1 OR_tmp196 (.Y(ttmp196),.A(N6871),.B(N6872));
OR2X1 OR_tmp197 (.Y(ttmp197),.A(N3210),.B(ttmp196));
OR2X1 OR_tmp198 (.Y(N7668),.A(N6870),.B(ttmp197));
OR2X1 OR_tmp199 (.Y(ttmp199),.A(N6886),.B(N6887));
OR2X1 OR_tmp200 (.Y(ttmp200),.A(N3228),.B(ttmp199));
OR2X1 OR_tmp201 (.Y(ttmp201),.A(N6884),.B(ttmp200));
OR2X1 OR_tmp202 (.Y(N7671),.A(N6885),.B(ttmp201));
NAND2X1 NAND2_2025 (.Y(N7744),.A(N3661),.B(N6968));
NAND2X1 NAND2_2026 (.Y(N7822),.A(N3664),.B(N7056));
OR2X1 OR_tmp203 (.Y(ttmp203),.A(N7061),.B(N7062));
OR2X1 OR_tmp204 (.Y(ttmp204),.A(N3361),.B(ttmp203));
OR2X1 OR_tmp205 (.Y(N7825),.A(N7060),.B(ttmp204));
OR2X1 OR_tmp206 (.Y(ttmp206),.A(N7066),.B(N7067));
OR2X1 OR_tmp207 (.Y(ttmp207),.A(N3365),.B(ttmp206));
OR2X1 OR_tmp208 (.Y(ttmp208),.A(N7064),.B(ttmp207));
OR2X1 OR_tmp209 (.Y(N7826),.A(N7065),.B(ttmp208));
OR2X1 OR_tmp210 (.Y(ttmp210),.A(N7105),.B(N7106));
OR2X1 OR_tmp211 (.Y(ttmp211),.A(N3370),.B(ttmp210));
OR2X1 OR_tmp212 (.Y(ttmp212),.A(N7103),.B(ttmp211));
OR2X1 OR_tmp213 (.Y(N7852),.A(N7104),.B(ttmp212));
OR2X1 OR_tmp214 (.Y(ttmp214),.A(N6778),.B(N6779));
OR2X1 OR_tmp215 (.Y(ttmp215),.A(N3101),.B(ttmp214));
OR2X1 OR_tmp216 (.Y(N8114),.A(N6777),.B(ttmp215));
OR2X1 OR_tmp217 (.Y(ttmp217),.A(N6772),.B(N6773));
OR2X1 OR_tmp218 (.Y(ttmp218),.A(N3097),.B(ttmp217));
OR2X1 OR_tmp219 (.Y(ttmp219),.A(N6770),.B(ttmp218));
OR2X1 OR_tmp220 (.Y(N8117),.A(N6771),.B(ttmp219));
OR2X1 OR_tmp221 (.Y(ttmp221),.A(N6780),.B(N6781));
NOR2X1 NOR_tmp222 (.Y(N8131),.A(N3101),.B(ttmp221));
OR2X1 OR_tmp223 (.Y(ttmp223),.A(N6775),.B(N6776));
OR2X1 OR_tmp224 (.Y(ttmp224),.A(N3097),.B(ttmp223));
NOR2X1 NOR_tmp225 (.Y(N8134),.A(N6774),.B(ttmp224));
NAND2X1 NAND2_2034 (.Y(N8144),.A(N6199),.B(N7477));
NAND2X1 NAND2_2035 (.Y(N8145),.A(N6196),.B(N7478));
OR2X1 OR_tmp226 (.Y(ttmp226),.A(N6840),.B(N6841));
OR2X1 OR_tmp227 (.Y(ttmp227),.A(N3169),.B(ttmp226));
OR2X1 OR_tmp228 (.Y(N8146),.A(N6839),.B(ttmp227));
OR2X1 OR_tmp229 (.Y(ttmp229),.A(N6842),.B(N6843));
NOR2X1 NOR_tmp230 (.Y(N8156),.A(N3169),.B(ttmp229));
OR2X1 OR_tmp231 (.Y(ttmp231),.A(N6860),.B(N6861));
OR2X1 OR_tmp232 (.Y(ttmp232),.A(N3189),.B(ttmp231));
OR2X1 OR_tmp233 (.Y(N8166),.A(N6859),.B(ttmp232));
OR2X1 OR_tmp234 (.Y(ttmp234),.A(N6854),.B(N6855));
OR2X1 OR_tmp235 (.Y(ttmp235),.A(N3185),.B(ttmp234));
OR2X1 OR_tmp236 (.Y(ttmp236),.A(N6852),.B(ttmp235));
OR2X1 OR_tmp237 (.Y(N8169),.A(N6853),.B(ttmp236));
OR2X1 OR_tmp238 (.Y(ttmp238),.A(N6862),.B(N6863));
NOR2X1 NOR_tmp239 (.Y(N8183),.A(N3189),.B(ttmp238));
OR2X1 OR_tmp240 (.Y(ttmp240),.A(N6857),.B(N6858));
OR2X1 OR_tmp241 (.Y(ttmp241),.A(N3185),.B(ttmp240));
NOR2X1 NOR_tmp242 (.Y(N8186),.A(N6856),.B(ttmp241));
OR2X1 OR_tmp243 (.Y(ttmp243),.A(N6874),.B(N6875));
OR2X1 OR_tmp244 (.Y(ttmp244),.A(N3211),.B(ttmp243));
OR2X1 OR_tmp245 (.Y(N8196),.A(N6873),.B(ttmp244));
OR2X1 OR_tmp246 (.Y(ttmp246),.A(N6876),.B(N6877));
NOR2X1 NOR_tmp247 (.Y(N8200),.A(N3211),.B(ttmp246));
OR2X1 OR_tmp248 (.Y(ttmp248),.A(N6878),.B(N6879));
OR2X1 OR_tmp249 (.Y(N8204),.A(N3215),.B(ttmp248));
NOR2X1 NOR2_2045 (.Y(N8208),.A(N3215),.B(N6880));
NAND2X1 NAND2_2046 (.Y(N8216),.A(N6252),.B(N7556));
NAND2X1 NAND2_2047 (.Y(N8217),.A(N6249),.B(N7557));
NAND2X1 NAND2_2048 (.Y(N8218),.A(N6246),.B(N7558));
NAND2X1 NAND2_2049 (.Y(N8219),.A(N6243),.B(N7559));
NAND2X1 NAND2_2050 (.Y(N8232),.A(N6266),.B(N7580));
NAND2X1 NAND2_2051 (.Y(N8233),.A(N6263),.B(N7581));
INVX1 NOT1_2052 (.Y(N8242),.A(N7411));
INVX1 NOT1_2053 (.Y(N8243),.A(N7414));
INVX1 NOT1_2054 (.Y(N8244),.A(N7417));
INVX1 NOT1_2055 (.Y(N8245),.A(N7420));
INVX1 NOT1_2056 (.Y(N8246),.A(N7423));
INVX1 NOT1_2057 (.Y(N8247),.A(N7426));
INVX1 NOT1_2058 (.Y(N8248),.A(N7429));
INVX1 NOT1_2059 (.Y(N8249),.A(N7432));
INVX1 NOT1_2060 (.Y(N8250),.A(N7435));
INVX1 NOT1_2061 (.Y(N8251),.A(N7438));
INVX1 NOT1_2062 (.Y(N8252),.A(N7136));
INVX1 NOT1_2063 (.Y(N8253),.A(N6923));
INVX1 NOT1_2064 (.Y(N8254),.A(N6762));
INVX1 NOT1_2065 (.Y(N8260),.A(N7459));
INVX1 NOT1_2066 (.Y(N8261),.A(N7462));
AND2X1 AND2_2067 (.Y(N8262),.A(N3122),.B(N6762));
AND2X1 AND2_2068 (.Y(N8269),.A(N3155),.B(N6784));
INVX1 NOT1_2069 (.Y(N8274),.A(N6815));
INVX1 NOT1_2070 (.Y(N8275),.A(N6818));
INVX1 NOT1_2071 (.Y(N8276),.A(N6821));
INVX1 NOT1_2072 (.Y(N8277),.A(N6824));
INVX1 NOT1_2073 (.Y(N8278),.A(N6827));
INVX1 NOT1_2074 (.Y(N8279),.A(N6830));
AND2X1 AND_tmp250 (.Y(ttmp250),.A(N5736),.B(N6815));
AND2X1 AND_tmp251 (.Y(N8280),.A(N5740),.B(ttmp250));
AND2X1 AND_tmp252 (.Y(ttmp252),.A(N6797),.B(N6818));
AND2X1 AND_tmp253 (.Y(N8281),.A(N6800),.B(ttmp252));
AND2X1 AND_tmp254 (.Y(ttmp254),.A(N5747),.B(N6821));
AND2X1 AND_tmp255 (.Y(N8282),.A(N5751),.B(ttmp254));
AND2X1 AND_tmp256 (.Y(ttmp256),.A(N6803),.B(N6824));
AND2X1 AND_tmp257 (.Y(N8283),.A(N6806),.B(ttmp256));
AND2X1 AND_tmp258 (.Y(ttmp258),.A(N5758),.B(N6827));
AND2X1 AND_tmp259 (.Y(N8284),.A(N5762),.B(ttmp258));
AND2X1 AND_tmp260 (.Y(ttmp260),.A(N6809),.B(N6830));
AND2X1 AND_tmp261 (.Y(N8285),.A(N6812),.B(ttmp260));
INVX1 NOT1_2081 (.Y(N8288),.A(N6845));
INVX1 NOT1_2082 (.Y(N8294),.A(N7488));
INVX1 NOT1_2083 (.Y(N8295),.A(N7500));
INVX1 NOT1_2084 (.Y(N8296),.A(N7515));
INVX1 NOT1_2085 (.Y(N8297),.A(N7518));
AND2X1 AND2_2086 (.Y(N8298),.A(N6833),.B(N6845));
AND2X1 AND2_2087 (.Y(N8307),.A(N6867),.B(N6881));
INVX1 NOT1_2088 (.Y(N8315),.A(N7533));
INVX1 NOT1_2089 (.Y(N8317),.A(N7536));
INVX1 NOT1_2090 (.Y(N8319),.A(N7539));
INVX1 NOT1_2091 (.Y(N8321),.A(N7542));
NAND2X1 NAND2_2092 (.Y(N8322),.A(N7545),.B(N4543));
INVX1 NOT1_2093 (.Y(N8323),.A(N7545));
NAND2X1 NAND2_2094 (.Y(N8324),.A(N7548),.B(N5943));
INVX1 NOT1_2095 (.Y(N8325),.A(N7548));
NAND2X1 NAND2_2096 (.Y(N8326),.A(N6967),.B(N7744));
AND2X1 AND_tmp262 (.Y(ttmp262),.A(N6912),.B(N6894));
AND2X1 AND_tmp263 (.Y(ttmp263),.A(N6901),.B(ttmp262));
AND2X1 AND_tmp264 (.Y(N8333),.A(N6923),.B(ttmp263));
AND2X1 AND2_2098 (.Y(N8337),.A(N6894),.B(N4545));
AND2X1 AND_tmp265 (.Y(ttmp265),.A(N6894),.B(N4549));
AND2X1 AND_tmp266 (.Y(N8338),.A(N6901),.B(ttmp265));
AND2X1 AND_tmp267 (.Y(ttmp267),.A(N4555),.B(N6901));
AND2X1 AND_tmp268 (.Y(ttmp268),.A(N6912),.B(ttmp267));
AND2X1 AND_tmp269 (.Y(N8339),.A(N6894),.B(ttmp268));
AND2X1 AND2_2101 (.Y(N8340),.A(N6901),.B(N4549));
AND2X1 AND_tmp270 (.Y(ttmp270),.A(N4555),.B(N6901));
AND2X1 AND_tmp271 (.Y(N8341),.A(N6912),.B(ttmp270));
AND2X1 AND_tmp272 (.Y(ttmp272),.A(N6912),.B(N6901));
AND2X1 AND_tmp273 (.Y(N8342),.A(N6923),.B(ttmp272));
AND2X1 AND2_2104 (.Y(N8343),.A(N6901),.B(N4549));
AND2X1 AND_tmp274 (.Y(ttmp274),.A(N6912),.B(N6901));
AND2X1 AND_tmp275 (.Y(N8344),.A(N4555),.B(ttmp274));
AND2X1 AND2_2106 (.Y(N8345),.A(N6912),.B(N4555));
AND2X1 AND2_2107 (.Y(N8346),.A(N6923),.B(N6912));
AND2X1 AND2_2108 (.Y(N8347),.A(N6912),.B(N4555));
AND2X1 AND2_2109 (.Y(N8348),.A(N6929),.B(N4563));
AND2X1 AND_tmp276 (.Y(ttmp276),.A(N6929),.B(N4566));
AND2X1 AND_tmp277 (.Y(N8349),.A(N6936),.B(ttmp276));
AND2X1 AND_tmp278 (.Y(ttmp278),.A(N4570),.B(N6936));
AND2X1 AND_tmp279 (.Y(ttmp279),.A(N6946),.B(ttmp278));
AND2X1 AND_tmp280 (.Y(N8350),.A(N6929),.B(ttmp279));
AND2X1 AND_tmp281 (.Y(ttmp281),.A(N5960),.B(N6936));
AND2X1 AND_tmp282 (.Y(ttmp282),.A(N6957),.B(ttmp281));
AND2X1 AND_tmp283 (.Y(ttmp283),.A(N6946),.B(ttmp282));
AND2X1 AND_tmp284 (.Y(N8351),.A(N6929),.B(ttmp283));
AND2X1 AND2_2113 (.Y(N8352),.A(N6936),.B(N4566));
AND2X1 AND_tmp285 (.Y(ttmp285),.A(N4570),.B(N6936));
AND2X1 AND_tmp286 (.Y(N8353),.A(N6946),.B(ttmp285));
AND2X1 AND_tmp287 (.Y(ttmp287),.A(N5960),.B(N6936));
AND2X1 AND_tmp288 (.Y(ttmp288),.A(N6957),.B(ttmp287));
AND2X1 AND_tmp289 (.Y(N8354),.A(N6946),.B(ttmp288));
AND2X1 AND2_2116 (.Y(N8355),.A(N4570),.B(N6946));
AND2X1 AND_tmp290 (.Y(ttmp290),.A(N6946),.B(N5960));
AND2X1 AND_tmp291 (.Y(N8356),.A(N6957),.B(ttmp290));
AND2X1 AND2_2118 (.Y(N8357),.A(N6957),.B(N5960));
NAND2X1 NAND2_2119 (.Y(N8358),.A(N7055),.B(N7822));
AND2X1 AND_tmp292 (.Y(ttmp292),.A(N6977),.B(N6970));
AND2X1 AND_tmp293 (.Y(ttmp293),.A(N7049),.B(ttmp292));
AND2X1 AND_tmp294 (.Y(N8365),.A(N6988),.B(ttmp293));
AND2X1 AND2_2121 (.Y(N8369),.A(N6970),.B(N4577));
AND2X1 AND_tmp295 (.Y(ttmp295),.A(N6970),.B(N4581));
AND2X1 AND_tmp296 (.Y(N8370),.A(N6977),.B(ttmp295));
AND2X1 AND_tmp297 (.Y(ttmp297),.A(N4586),.B(N6977));
AND2X1 AND_tmp298 (.Y(ttmp298),.A(N6988),.B(ttmp297));
AND2X1 AND_tmp299 (.Y(N8371),.A(N6970),.B(ttmp298));
AND2X1 AND2_2124 (.Y(N8372),.A(N6977),.B(N4581));
AND2X1 AND_tmp300 (.Y(ttmp300),.A(N4586),.B(N6977));
AND2X1 AND_tmp301 (.Y(N8373),.A(N6988),.B(ttmp300));
AND2X1 AND_tmp302 (.Y(ttmp302),.A(N6988),.B(N6977));
AND2X1 AND_tmp303 (.Y(N8374),.A(N7049),.B(ttmp302));
AND2X1 AND2_2127 (.Y(N8375),.A(N6977),.B(N4581));
AND2X1 AND_tmp304 (.Y(ttmp304),.A(N4586),.B(N6977));
AND2X1 AND_tmp305 (.Y(N8376),.A(N6988),.B(ttmp304));
AND2X1 AND2_2129 (.Y(N8377),.A(N6988),.B(N4586));
AND2X1 AND2_2130 (.Y(N8378),.A(N6998),.B(N4593));
AND2X1 AND_tmp306 (.Y(ttmp306),.A(N6998),.B(N4597));
AND2X1 AND_tmp307 (.Y(N8379),.A(N7006),.B(ttmp306));
AND2X1 AND_tmp308 (.Y(ttmp308),.A(N4603),.B(N7006));
AND2X1 AND_tmp309 (.Y(ttmp309),.A(N7020),.B(ttmp308));
AND2X1 AND_tmp310 (.Y(N8380),.A(N6998),.B(ttmp309));
AND2X1 AND_tmp311 (.Y(ttmp311),.A(N5981),.B(N7006));
AND2X1 AND_tmp312 (.Y(ttmp312),.A(N7036),.B(ttmp311));
AND2X1 AND_tmp313 (.Y(ttmp313),.A(N7020),.B(ttmp312));
AND2X1 AND_tmp314 (.Y(N8381),.A(N6998),.B(ttmp313));
AND2X1 AND2_2134 (.Y(N8382),.A(N7006),.B(N4597));
AND2X1 AND_tmp315 (.Y(ttmp315),.A(N4603),.B(N7006));
AND2X1 AND_tmp316 (.Y(N8383),.A(N7020),.B(ttmp315));
AND2X1 AND_tmp317 (.Y(ttmp317),.A(N5981),.B(N7006));
AND2X1 AND_tmp318 (.Y(ttmp318),.A(N7036),.B(ttmp317));
AND2X1 AND_tmp319 (.Y(N8384),.A(N7020),.B(ttmp318));
AND2X1 AND2_2137 (.Y(N8385),.A(N7006),.B(N4597));
AND2X1 AND_tmp320 (.Y(ttmp320),.A(N4603),.B(N7006));
AND2X1 AND_tmp321 (.Y(N8386),.A(N7020),.B(ttmp320));
AND2X1 AND_tmp322 (.Y(ttmp322),.A(N5981),.B(N7006));
AND2X1 AND_tmp323 (.Y(ttmp323),.A(N7036),.B(ttmp322));
AND2X1 AND_tmp324 (.Y(N8387),.A(N7020),.B(ttmp323));
AND2X1 AND2_2140 (.Y(N8388),.A(N7020),.B(N4603));
AND2X1 AND_tmp325 (.Y(ttmp325),.A(N7020),.B(N5981));
AND2X1 AND_tmp326 (.Y(N8389),.A(N7036),.B(ttmp325));
AND2X1 AND2_2142 (.Y(N8390),.A(N7020),.B(N4603));
AND2X1 AND_tmp327 (.Y(ttmp327),.A(N7020),.B(N5981));
AND2X1 AND_tmp328 (.Y(N8391),.A(N7036),.B(ttmp327));
AND2X1 AND2_2144 (.Y(N8392),.A(N7036),.B(N5981));
AND2X1 AND2_2145 (.Y(N8393),.A(N7049),.B(N6988));
AND2X1 AND2_2146 (.Y(N8394),.A(N7057),.B(N7063));
AND2X1 AND2_2147 (.Y(N8404),.A(N7057),.B(N7826));
AND2X1 AND_tmp329 (.Y(ttmp329),.A(N7073),.B(N7068));
AND2X1 AND_tmp330 (.Y(ttmp330),.A(N7098),.B(ttmp329));
AND2X1 AND_tmp331 (.Y(N8405),.A(N7077),.B(ttmp330));
AND2X1 AND2_2149 (.Y(N8409),.A(N7068),.B(N4632));
AND2X1 AND_tmp332 (.Y(ttmp332),.A(N7068),.B(N4634));
AND2X1 AND_tmp333 (.Y(N8410),.A(N7073),.B(ttmp332));
AND2X1 AND_tmp334 (.Y(ttmp334),.A(N4635),.B(N7073));
AND2X1 AND_tmp335 (.Y(ttmp335),.A(N7077),.B(ttmp334));
AND2X1 AND_tmp336 (.Y(N8411),.A(N7068),.B(ttmp335));
AND2X1 AND_tmp337 (.Y(ttmp337),.A(N7086),.B(N7080));
AND2X1 AND_tmp338 (.Y(ttmp338),.A(N7099),.B(ttmp337));
AND2X1 AND_tmp339 (.Y(ttmp339),.A(N7095),.B(ttmp338));
AND2X1 AND_tmp340 (.Y(N8412),.A(N7091),.B(ttmp339));
AND2X1 AND2_2153 (.Y(N8415),.A(N7080),.B(N4638));
AND2X1 AND_tmp341 (.Y(ttmp341),.A(N7080),.B(N4639));
AND2X1 AND_tmp342 (.Y(N8416),.A(N7086),.B(ttmp341));
AND2X1 AND_tmp343 (.Y(ttmp343),.A(N4640),.B(N7086));
AND2X1 AND_tmp344 (.Y(ttmp344),.A(N7091),.B(ttmp343));
AND2X1 AND_tmp345 (.Y(N8417),.A(N7080),.B(ttmp344));
AND2X1 AND_tmp346 (.Y(ttmp346),.A(N4641),.B(N7086));
AND2X1 AND_tmp347 (.Y(ttmp347),.A(N7095),.B(ttmp346));
AND2X1 AND_tmp348 (.Y(ttmp348),.A(N7091),.B(ttmp347));
AND2X1 AND_tmp349 (.Y(N8418),.A(N7080),.B(ttmp348));
AND2X1 AND2_2157 (.Y(N8421),.A(N3375),.B(N7100));
AND2X1 AND_tmp350 (.Y(ttmp350),.A(N7125),.B(N7107));
AND2X1 AND_tmp351 (.Y(ttmp351),.A(N7114),.B(ttmp350));
AND2X1 AND_tmp352 (.Y(N8430),.A(N7136),.B(ttmp351));
AND2X1 AND2_2159 (.Y(N8433),.A(N7107),.B(N4657));
AND2X1 AND_tmp353 (.Y(ttmp353),.A(N7107),.B(N4661));
AND2X1 AND_tmp354 (.Y(N8434),.A(N7114),.B(ttmp353));
AND2X1 AND_tmp355 (.Y(ttmp355),.A(N4667),.B(N7114));
AND2X1 AND_tmp356 (.Y(ttmp356),.A(N7125),.B(ttmp355));
AND2X1 AND_tmp357 (.Y(N8435),.A(N7107),.B(ttmp356));
AND2X1 AND2_2162 (.Y(N8436),.A(N7114),.B(N4661));
AND2X1 AND_tmp358 (.Y(ttmp358),.A(N4667),.B(N7114));
AND2X1 AND_tmp359 (.Y(N8437),.A(N7125),.B(ttmp358));
AND2X1 AND_tmp360 (.Y(ttmp360),.A(N7125),.B(N7114));
AND2X1 AND_tmp361 (.Y(N8438),.A(N7136),.B(ttmp360));
AND2X1 AND2_2165 (.Y(N8439),.A(N7114),.B(N4661));
AND2X1 AND_tmp362 (.Y(ttmp362),.A(N7125),.B(N7114));
AND2X1 AND_tmp363 (.Y(N8440),.A(N4667),.B(ttmp362));
AND2X1 AND2_2167 (.Y(N8441),.A(N7125),.B(N4667));
AND2X1 AND2_2168 (.Y(N8442),.A(N7136),.B(N7125));
AND2X1 AND2_2169 (.Y(N8443),.A(N7125),.B(N4667));
AND2X1 AND_tmp364 (.Y(ttmp364),.A(N7142),.B(N7170));
AND2X1 AND_tmp365 (.Y(ttmp365),.A(N7149),.B(ttmp364));
AND2X1 AND_tmp366 (.Y(ttmp366),.A(N7180),.B(ttmp365));
AND2X1 AND_tmp367 (.Y(N8444),.A(N7159),.B(ttmp366));
AND2X1 AND2_2171 (.Y(N8447),.A(N7142),.B(N4675));
AND2X1 AND_tmp368 (.Y(ttmp368),.A(N7142),.B(N4678));
AND2X1 AND_tmp369 (.Y(N8448),.A(N7149),.B(ttmp368));
AND2X1 AND_tmp370 (.Y(ttmp370),.A(N4682),.B(N7149));
AND2X1 AND_tmp371 (.Y(ttmp371),.A(N7159),.B(ttmp370));
AND2X1 AND_tmp372 (.Y(N8449),.A(N7142),.B(ttmp371));
AND2X1 AND_tmp373 (.Y(ttmp373),.A(N4687),.B(N7149));
AND2X1 AND_tmp374 (.Y(ttmp374),.A(N7170),.B(ttmp373));
AND2X1 AND_tmp375 (.Y(ttmp375),.A(N7159),.B(ttmp374));
AND2X1 AND_tmp376 (.Y(N8450),.A(N7142),.B(ttmp375));
AND2X1 AND2_2175 (.Y(N8451),.A(N7149),.B(N4678));
AND2X1 AND_tmp377 (.Y(ttmp377),.A(N4682),.B(N7149));
AND2X1 AND_tmp378 (.Y(N8452),.A(N7159),.B(ttmp377));
AND2X1 AND_tmp379 (.Y(ttmp379),.A(N4687),.B(N7149));
AND2X1 AND_tmp380 (.Y(ttmp380),.A(N7170),.B(ttmp379));
AND2X1 AND_tmp381 (.Y(N8453),.A(N7159),.B(ttmp380));
AND2X1 AND2_2178 (.Y(N8454),.A(N4682),.B(N7159));
AND2X1 AND_tmp382 (.Y(ttmp382),.A(N7159),.B(N4687));
AND2X1 AND_tmp383 (.Y(N8455),.A(N7170),.B(ttmp382));
AND2X1 AND2_2180 (.Y(N8456),.A(N7170),.B(N4687));
INVX1 NOT1_2181 (.Y(N8457),.A(N7194));
INVX1 NOT1_2182 (.Y(N8460),.A(N7198));
INVX1 NOT1_2183 (.Y(N8463),.A(N7205));
INVX1 NOT1_2184 (.Y(N8466),.A(N7209));
INVX1 NOT1_2185 (.Y(N8469),.A(N7216));
INVX1 NOT1_2186 (.Y(N8470),.A(N7219));
BUFX1 BUFF1_2187 (.Y(N8471),.A(N7202));
BUFX1 BUFF1_2188 (.Y(N8474),.A(N7202));
BUFX1 BUFF1_2189 (.Y(N8477),.A(N7213));
BUFX1 BUFF1_2190 (.Y(N8480),.A(N7213));
AND2X1 AND_tmp384 (.Y(ttmp384),.A(N6079),.B(N7216));
AND2X1 AND_tmp385 (.Y(N8483),.A(N6083),.B(ttmp384));
AND2X1 AND_tmp386 (.Y(ttmp386),.A(N7188),.B(N7219));
AND2X1 AND_tmp387 (.Y(N8484),.A(N7191),.B(ttmp386));
AND2X1 AND_tmp388 (.Y(ttmp388),.A(N7229),.B(N7222));
AND2X1 AND_tmp389 (.Y(ttmp389),.A(N7301),.B(ttmp388));
AND2X1 AND_tmp390 (.Y(N8485),.A(N7240),.B(ttmp389));
AND2X1 AND2_2194 (.Y(N8488),.A(N7222),.B(N4702));
AND2X1 AND_tmp391 (.Y(ttmp391),.A(N7222),.B(N4706));
AND2X1 AND_tmp392 (.Y(N8489),.A(N7229),.B(ttmp391));
AND2X1 AND_tmp393 (.Y(ttmp393),.A(N4711),.B(N7229));
AND2X1 AND_tmp394 (.Y(ttmp394),.A(N7240),.B(ttmp393));
AND2X1 AND_tmp395 (.Y(N8490),.A(N7222),.B(ttmp394));
AND2X1 AND2_2197 (.Y(N8491),.A(N7229),.B(N4706));
AND2X1 AND_tmp396 (.Y(ttmp396),.A(N4711),.B(N7229));
AND2X1 AND_tmp397 (.Y(N8492),.A(N7240),.B(ttmp396));
AND2X1 AND_tmp398 (.Y(ttmp398),.A(N7240),.B(N7229));
AND2X1 AND_tmp399 (.Y(N8493),.A(N7301),.B(ttmp398));
AND2X1 AND2_2200 (.Y(N8494),.A(N7229),.B(N4706));
AND2X1 AND_tmp400 (.Y(ttmp400),.A(N4711),.B(N7229));
AND2X1 AND_tmp401 (.Y(N8495),.A(N7240),.B(ttmp400));
AND2X1 AND2_2202 (.Y(N8496),.A(N7240),.B(N4711));
AND2X1 AND_tmp402 (.Y(ttmp402),.A(N7258),.B(N7250));
AND2X1 AND_tmp403 (.Y(ttmp403),.A(N7307),.B(ttmp402));
AND2X1 AND_tmp404 (.Y(ttmp404),.A(N7288),.B(ttmp403));
AND2X1 AND_tmp405 (.Y(N8497),.A(N7272),.B(ttmp404));
AND2X1 AND2_2204 (.Y(N8500),.A(N7250),.B(N4718));
AND2X1 AND_tmp406 (.Y(ttmp406),.A(N7250),.B(N4722));
AND2X1 AND_tmp407 (.Y(N8501),.A(N7258),.B(ttmp406));
AND2X1 AND_tmp408 (.Y(ttmp408),.A(N4728),.B(N7258));
AND2X1 AND_tmp409 (.Y(ttmp409),.A(N7272),.B(ttmp408));
AND2X1 AND_tmp410 (.Y(N8502),.A(N7250),.B(ttmp409));
AND2X1 AND_tmp411 (.Y(ttmp411),.A(N4735),.B(N7258));
AND2X1 AND_tmp412 (.Y(ttmp412),.A(N7288),.B(ttmp411));
AND2X1 AND_tmp413 (.Y(ttmp413),.A(N7272),.B(ttmp412));
AND2X1 AND_tmp414 (.Y(N8503),.A(N7250),.B(ttmp413));
AND2X1 AND2_2208 (.Y(N8504),.A(N7258),.B(N4722));
AND2X1 AND_tmp415 (.Y(ttmp415),.A(N4728),.B(N7258));
AND2X1 AND_tmp416 (.Y(N8505),.A(N7272),.B(ttmp415));
AND2X1 AND_tmp417 (.Y(ttmp417),.A(N4735),.B(N7258));
AND2X1 AND_tmp418 (.Y(ttmp418),.A(N7288),.B(ttmp417));
AND2X1 AND_tmp419 (.Y(N8506),.A(N7272),.B(ttmp418));
AND2X1 AND_tmp420 (.Y(ttmp420),.A(N7258),.B(N7288));
AND2X1 AND_tmp421 (.Y(ttmp421),.A(N7307),.B(ttmp420));
AND2X1 AND_tmp422 (.Y(N8507),.A(N7272),.B(ttmp421));
AND2X1 AND2_2212 (.Y(N8508),.A(N7258),.B(N4722));
AND2X1 AND_tmp423 (.Y(ttmp423),.A(N4728),.B(N7258));
AND2X1 AND_tmp424 (.Y(N8509),.A(N7272),.B(ttmp423));
AND2X1 AND_tmp425 (.Y(ttmp425),.A(N4735),.B(N7258));
AND2X1 AND_tmp426 (.Y(ttmp426),.A(N7288),.B(ttmp425));
AND2X1 AND_tmp427 (.Y(N8510),.A(N7272),.B(ttmp426));
AND2X1 AND2_2215 (.Y(N8511),.A(N7272),.B(N4728));
AND2X1 AND_tmp428 (.Y(ttmp428),.A(N7272),.B(N4735));
AND2X1 AND_tmp429 (.Y(N8512),.A(N7288),.B(ttmp428));
AND2X1 AND_tmp430 (.Y(ttmp430),.A(N7272),.B(N7288));
AND2X1 AND_tmp431 (.Y(N8513),.A(N7307),.B(ttmp430));
AND2X1 AND2_2218 (.Y(N8514),.A(N7272),.B(N4728));
AND2X1 AND_tmp432 (.Y(ttmp432),.A(N7272),.B(N4735));
AND2X1 AND_tmp433 (.Y(N8515),.A(N7288),.B(ttmp432));
AND2X1 AND2_2220 (.Y(N8516),.A(N7288),.B(N4735));
AND2X1 AND2_2221 (.Y(N8517),.A(N7301),.B(N7240));
AND2X1 AND2_2222 (.Y(N8518),.A(N7307),.B(N7288));
INVX1 NOT1_2223 (.Y(N8519),.A(N7314));
INVX1 NOT1_2224 (.Y(N8522),.A(N7318));
BUFX1 BUFF1_2225 (.Y(N8525),.A(N7322));
BUFX1 BUFF1_2226 (.Y(N8528),.A(N7322));
BUFX1 BUFF1_2227 (.Y(N8531),.A(N7331));
BUFX1 BUFF1_2228 (.Y(N8534),.A(N7331));
INVX1 NOT1_2229 (.Y(N8537),.A(N7340));
INVX1 NOT1_2230 (.Y(N8538),.A(N7343));
AND2X1 AND_tmp434 (.Y(ttmp434),.A(N6137),.B(N7340));
AND2X1 AND_tmp435 (.Y(N8539),.A(N6141),.B(ttmp434));
AND2X1 AND_tmp436 (.Y(ttmp436),.A(N7334),.B(N7343));
AND2X1 AND_tmp437 (.Y(N8540),.A(N7337),.B(ttmp436));
AND2X1 AND_tmp438 (.Y(ttmp438),.A(N7351),.B(N7346));
AND2X1 AND_tmp439 (.Y(ttmp439),.A(N7376),.B(ttmp438));
AND2X1 AND_tmp440 (.Y(N8541),.A(N7355),.B(ttmp439));
AND2X1 AND2_2234 (.Y(N8545),.A(N7346),.B(N4757));
AND2X1 AND_tmp441 (.Y(ttmp441),.A(N7346),.B(N4758));
AND2X1 AND_tmp442 (.Y(N8546),.A(N7351),.B(ttmp441));
AND2X1 AND_tmp443 (.Y(ttmp443),.A(N4759),.B(N7351));
AND2X1 AND_tmp444 (.Y(ttmp444),.A(N7355),.B(ttmp443));
AND2X1 AND_tmp445 (.Y(N8547),.A(N7346),.B(ttmp444));
AND2X1 AND_tmp446 (.Y(ttmp446),.A(N7364),.B(N7358));
AND2X1 AND_tmp447 (.Y(ttmp447),.A(N7377),.B(ttmp446));
AND2X1 AND_tmp448 (.Y(ttmp448),.A(N7373),.B(ttmp447));
AND2X1 AND_tmp449 (.Y(N8548),.A(N7369),.B(ttmp448));
AND2X1 AND2_2238 (.Y(N8551),.A(N7358),.B(N4762));
AND2X1 AND_tmp450 (.Y(ttmp450),.A(N7358),.B(N4764));
AND2X1 AND_tmp451 (.Y(N8552),.A(N7364),.B(ttmp450));
AND2X1 AND_tmp452 (.Y(ttmp452),.A(N4766),.B(N7364));
AND2X1 AND_tmp453 (.Y(ttmp453),.A(N7369),.B(ttmp452));
AND2X1 AND_tmp454 (.Y(N8553),.A(N7358),.B(ttmp453));
AND2X1 AND_tmp455 (.Y(ttmp455),.A(N4767),.B(N7364));
AND2X1 AND_tmp456 (.Y(ttmp456),.A(N7373),.B(ttmp455));
AND2X1 AND_tmp457 (.Y(ttmp457),.A(N7369),.B(ttmp456));
AND2X1 AND_tmp458 (.Y(N8554),.A(N7358),.B(ttmp457));
INVX1 NOT1_2242 (.Y(N8555),.A(N7387));
INVX1 NOT1_2243 (.Y(N8558),.A(N7394));
INVX1 NOT1_2244 (.Y(N8561),.A(N7398));
INVX1 NOT1_2245 (.Y(N8564),.A(N7405));
INVX1 NOT1_2246 (.Y(N8565),.A(N7408));
BUFX1 BUFF1_2247 (.Y(N8566),.A(N7391));
BUFX1 BUFF1_2248 (.Y(N8569),.A(N7391));
BUFX1 BUFF1_2249 (.Y(N8572),.A(N7402));
BUFX1 BUFF1_2250 (.Y(N8575),.A(N7402));
AND2X1 AND_tmp459 (.Y(ttmp459),.A(N6166),.B(N7405));
AND2X1 AND_tmp460 (.Y(N8578),.A(N6170),.B(ttmp459));
AND2X1 AND_tmp461 (.Y(ttmp461),.A(N7378),.B(N7408));
AND2X1 AND_tmp462 (.Y(N8579),.A(N7381),.B(ttmp461));
BUFX1 BUFF1_2253 (.Y(N8580),.A(N7180));
BUFX1 BUFF1_2254 (.Y(N8583),.A(N7142));
BUFX1 BUFF1_2255 (.Y(N8586),.A(N7149));
BUFX1 BUFF1_2256 (.Y(N8589),.A(N7159));
BUFX1 BUFF1_2257 (.Y(N8592),.A(N7170));
BUFX1 BUFF1_2258 (.Y(N8595),.A(N6929));
BUFX1 BUFF1_2259 (.Y(N8598),.A(N6936));
BUFX1 BUFF1_2260 (.Y(N8601),.A(N6946));
BUFX1 BUFF1_2261 (.Y(N8604),.A(N6957));
INVX1 NOT1_2262 (.Y(N8607),.A(N7441));
NAND2X1 NAND2_2263 (.Y(N8608),.A(N7441),.B(N5469));
INVX1 NOT1_2264 (.Y(N8609),.A(N7444));
NAND2X1 NAND2_2265 (.Y(N8610),.A(N7444),.B(N4793));
INVX1 NOT1_2266 (.Y(N8615),.A(N7447));
INVX1 NOT1_2267 (.Y(N8616),.A(N7450));
INVX1 NOT1_2268 (.Y(N8617),.A(N7453));
INVX1 NOT1_2269 (.Y(N8618),.A(N7456));
INVX1 NOT1_2270 (.Y(N8619),.A(N7474));
INVX1 NOT1_2271 (.Y(N8624),.A(N7465));
INVX1 NOT1_2272 (.Y(N8625),.A(N7468));
INVX1 NOT1_2273 (.Y(N8626),.A(N7471));
NAND2X1 NAND2_2274 (.Y(N8627),.A(N8144),.B(N8145));
INVX1 NOT1_2275 (.Y(N8632),.A(N7479));
INVX1 NOT1_2276 (.Y(N8633),.A(N7482));
INVX1 NOT1_2277 (.Y(N8634),.A(N7485));
INVX1 NOT1_2278 (.Y(N8637),.A(N7491));
INVX1 NOT1_2279 (.Y(N8638),.A(N7494));
INVX1 NOT1_2280 (.Y(N8639),.A(N7497));
INVX1 NOT1_2281 (.Y(N8644),.A(N7503));
INVX1 NOT1_2282 (.Y(N8645),.A(N7506));
INVX1 NOT1_2283 (.Y(N8646),.A(N7509));
INVX1 NOT1_2284 (.Y(N8647),.A(N7512));
INVX1 NOT1_2285 (.Y(N8648),.A(N7530));
INVX1 NOT1_2286 (.Y(N8653),.A(N7521));
INVX1 NOT1_2287 (.Y(N8654),.A(N7524));
INVX1 NOT1_2288 (.Y(N8655),.A(N7527));
BUFX1 BUFF1_2289 (.Y(N8660),.A(N6894));
BUFX1 BUFF1_2290 (.Y(N8663),.A(N6894));
BUFX1 BUFF1_2291 (.Y(N8666),.A(N6901));
BUFX1 BUFF1_2292 (.Y(N8669),.A(N6901));
BUFX1 BUFF1_2293 (.Y(N8672),.A(N6912));
BUFX1 BUFF1_2294 (.Y(N8675),.A(N6912));
BUFX1 BUFF1_2295 (.Y(N8678),.A(N7049));
BUFX1 BUFF1_2296 (.Y(N8681),.A(N6988));
BUFX1 BUFF1_2297 (.Y(N8684),.A(N6970));
BUFX1 BUFF1_2298 (.Y(N8687),.A(N6977));
BUFX1 BUFF1_2299 (.Y(N8690),.A(N7049));
BUFX1 BUFF1_2300 (.Y(N8693),.A(N6988));
BUFX1 BUFF1_2301 (.Y(N8696),.A(N6970));
BUFX1 BUFF1_2302 (.Y(N8699),.A(N6977));
BUFX1 BUFF1_2303 (.Y(N8702),.A(N7036));
BUFX1 BUFF1_2304 (.Y(N8705),.A(N6998));
BUFX1 BUFF1_2305 (.Y(N8708),.A(N7020));
BUFX1 BUFF1_2306 (.Y(N8711),.A(N7006));
BUFX1 BUFF1_2307 (.Y(N8714),.A(N7006));
INVX1 NOT1_2308 (.Y(N8717),.A(N7553));
BUFX1 BUFF1_2309 (.Y(N8718),.A(N7036));
BUFX1 BUFF1_2310 (.Y(N8721),.A(N6998));
BUFX1 BUFF1_2311 (.Y(N8724),.A(N7020));
NAND2X1 NAND2_2312 (.Y(N8727),.A(N8216),.B(N8217));
NAND2X1 NAND2_2313 (.Y(N8730),.A(N8218),.B(N8219));
INVX1 NOT1_2314 (.Y(N8733),.A(N7574));
INVX1 NOT1_2315 (.Y(N8734),.A(N7577));
BUFX1 BUFF1_2316 (.Y(N8735),.A(N7107));
BUFX1 BUFF1_2317 (.Y(N8738),.A(N7107));
BUFX1 BUFF1_2318 (.Y(N8741),.A(N7114));
BUFX1 BUFF1_2319 (.Y(N8744),.A(N7114));
BUFX1 BUFF1_2320 (.Y(N8747),.A(N7125));
BUFX1 BUFF1_2321 (.Y(N8750),.A(N7125));
INVX1 NOT1_2322 (.Y(N8753),.A(N7560));
INVX1 NOT1_2323 (.Y(N8754),.A(N7563));
INVX1 NOT1_2324 (.Y(N8755),.A(N7566));
INVX1 NOT1_2325 (.Y(N8756),.A(N7569));
BUFX1 BUFF1_2326 (.Y(N8757),.A(N7301));
BUFX1 BUFF1_2327 (.Y(N8760),.A(N7240));
BUFX1 BUFF1_2328 (.Y(N8763),.A(N7222));
BUFX1 BUFF1_2329 (.Y(N8766),.A(N7229));
BUFX1 BUFF1_2330 (.Y(N8769),.A(N7301));
BUFX1 BUFF1_2331 (.Y(N8772),.A(N7240));
BUFX1 BUFF1_2332 (.Y(N8775),.A(N7222));
BUFX1 BUFF1_2333 (.Y(N8778),.A(N7229));
BUFX1 BUFF1_2334 (.Y(N8781),.A(N7307));
BUFX1 BUFF1_2335 (.Y(N8784),.A(N7288));
BUFX1 BUFF1_2336 (.Y(N8787),.A(N7250));
BUFX1 BUFF1_2337 (.Y(N8790),.A(N7272));
BUFX1 BUFF1_2338 (.Y(N8793),.A(N7258));
BUFX1 BUFF1_2339 (.Y(N8796),.A(N7258));
BUFX1 BUFF1_2340 (.Y(N8799),.A(N7307));
BUFX1 BUFF1_2341 (.Y(N8802),.A(N7288));
BUFX1 BUFF1_2342 (.Y(N8805),.A(N7250));
BUFX1 BUFF1_2343 (.Y(N8808),.A(N7272));
NAND2X1 NAND2_2344 (.Y(N8811),.A(N8232),.B(N8233));
INVX1 NOT1_2345 (.Y(N8814),.A(N7588));
INVX1 NOT1_2346 (.Y(N8815),.A(N7591));
INVX1 NOT1_2347 (.Y(N8816),.A(N7582));
INVX1 NOT1_2348 (.Y(N8817),.A(N7585));
AND2X1 AND2_2349 (.Y(N8818),.A(N7620),.B(N3155));
AND2X1 AND2_2350 (.Y(N8840),.A(N3122),.B(N7609));
INVX1 NOT1_2351 (.Y(N8857),.A(N7609));
AND2X1 AND_tmp463 (.Y(ttmp463),.A(N5740),.B(N8274));
AND2X1 AND_tmp464 (.Y(N8861),.A(N6797),.B(ttmp463));
AND2X1 AND_tmp465 (.Y(ttmp465),.A(N6800),.B(N8275));
AND2X1 AND_tmp466 (.Y(N8862),.A(N5736),.B(ttmp465));
AND2X1 AND_tmp467 (.Y(ttmp467),.A(N5751),.B(N8276));
AND2X1 AND_tmp468 (.Y(N8863),.A(N6803),.B(ttmp467));
AND2X1 AND_tmp469 (.Y(ttmp469),.A(N6806),.B(N8277));
AND2X1 AND_tmp470 (.Y(N8864),.A(N5747),.B(ttmp469));
AND2X1 AND_tmp471 (.Y(ttmp471),.A(N5762),.B(N8278));
AND2X1 AND_tmp472 (.Y(N8865),.A(N6809),.B(ttmp471));
AND2X1 AND_tmp473 (.Y(ttmp473),.A(N6812),.B(N8279));
AND2X1 AND_tmp474 (.Y(N8866),.A(N5758),.B(ttmp473));
INVX1 NOT1_2358 (.Y(N8871),.A(N7655));
AND2X1 AND2_2359 (.Y(N8874),.A(N6833),.B(N7655));
AND2X1 AND2_2360 (.Y(N8878),.A(N7671),.B(N6867));
INVX1 NOT1_2361 (.Y(N8879),.A(N8196));
NAND2X1 NAND2_2362 (.Y(N8880),.A(N8196),.B(N8315));
INVX1 NOT1_2363 (.Y(N8881),.A(N8200));
NAND2X1 NAND2_2364 (.Y(N8882),.A(N8200),.B(N8317));
INVX1 NOT1_2365 (.Y(N8883),.A(N8204));
NAND2X1 NAND2_2366 (.Y(N8884),.A(N8204),.B(N8319));
INVX1 NOT1_2367 (.Y(N8885),.A(N8208));
NAND2X1 NAND2_2368 (.Y(N8886),.A(N8208),.B(N8321));
NAND2X1 NAND2_2369 (.Y(N8887),.A(N3658),.B(N8323));
NAND2X1 NAND2_2370 (.Y(N8888),.A(N4817),.B(N8325));
OR2X1 OR_tmp475 (.Y(ttmp475),.A(N8338),.B(N8339));
OR2X1 OR_tmp476 (.Y(ttmp476),.A(N4544),.B(ttmp475));
OR2X1 OR_tmp477 (.Y(N8898),.A(N8337),.B(ttmp476));
OR2X1 OR_tmp478 (.Y(ttmp478),.A(N8350),.B(N8351));
OR2X1 OR_tmp479 (.Y(ttmp479),.A(N4562),.B(ttmp478));
OR2X1 OR_tmp480 (.Y(ttmp480),.A(N8348),.B(ttmp479));
OR2X1 OR_tmp481 (.Y(N8902),.A(N8349),.B(ttmp480));
OR2X1 OR_tmp482 (.Y(ttmp482),.A(N8370),.B(N8371));
OR2X1 OR_tmp483 (.Y(ttmp483),.A(N4576),.B(ttmp482));
OR2X1 OR_tmp484 (.Y(N8920),.A(N8369),.B(ttmp483));
OR2X1 OR2_2374 (.Y(N8924),.A(N4581),.B(N8377));
OR2X1 OR_tmp485 (.Y(ttmp485),.A(N8380),.B(N8381));
OR2X1 OR_tmp486 (.Y(ttmp486),.A(N4592),.B(ttmp485));
OR2X1 OR_tmp487 (.Y(ttmp487),.A(N8378),.B(ttmp486));
OR2X1 OR_tmp488 (.Y(N8927),.A(N8379),.B(ttmp487));
OR2X1 OR2_2376 (.Y(N8931),.A(N4603),.B(N8392));
OR2X1 OR2_2377 (.Y(N8943),.A(N7825),.B(N8404));
OR2X1 OR_tmp489 (.Y(ttmp489),.A(N8410),.B(N8411));
OR2X1 OR_tmp490 (.Y(ttmp490),.A(N4630),.B(ttmp489));
OR2X1 OR_tmp491 (.Y(N8950),.A(N8409),.B(ttmp490));
OR2X1 OR_tmp492 (.Y(ttmp492),.A(N8417),.B(N8418));
OR2X1 OR_tmp493 (.Y(ttmp493),.A(N4637),.B(ttmp492));
OR2X1 OR_tmp494 (.Y(ttmp494),.A(N8415),.B(ttmp493));
OR2X1 OR_tmp495 (.Y(N8956),.A(N8416),.B(ttmp494));
INVX1 NOT1_2380 (.Y(N8959),.A(N7852));
AND2X1 AND2_2381 (.Y(N8960),.A(N3375),.B(N7852));
OR2X1 OR_tmp496 (.Y(ttmp496),.A(N8434),.B(N8435));
OR2X1 OR_tmp497 (.Y(ttmp497),.A(N4656),.B(ttmp496));
OR2X1 OR_tmp498 (.Y(N8963),.A(N8433),.B(ttmp497));
OR2X1 OR_tmp499 (.Y(ttmp499),.A(N8449),.B(N8450));
OR2X1 OR_tmp500 (.Y(ttmp500),.A(N4674),.B(ttmp499));
OR2X1 OR_tmp501 (.Y(ttmp501),.A(N8447),.B(ttmp500));
OR2X1 OR_tmp502 (.Y(N8966),.A(N8448),.B(ttmp501));
AND2X1 AND_tmp503 (.Y(ttmp503),.A(N6083),.B(N8469));
AND2X1 AND_tmp504 (.Y(N8991),.A(N7188),.B(ttmp503));
AND2X1 AND_tmp505 (.Y(ttmp505),.A(N7191),.B(N8470));
AND2X1 AND_tmp506 (.Y(N8992),.A(N6079),.B(ttmp505));
OR2X1 OR_tmp507 (.Y(ttmp507),.A(N8489),.B(N8490));
OR2X1 OR_tmp508 (.Y(ttmp508),.A(N4701),.B(ttmp507));
OR2X1 OR_tmp509 (.Y(N8995),.A(N8488),.B(ttmp508));
OR2X1 OR2_2387 (.Y(N8996),.A(N4706),.B(N8496));
OR2X1 OR_tmp510 (.Y(ttmp510),.A(N8502),.B(N8503));
OR2X1 OR_tmp511 (.Y(ttmp511),.A(N4717),.B(ttmp510));
OR2X1 OR_tmp512 (.Y(ttmp512),.A(N8500),.B(ttmp511));
OR2X1 OR_tmp513 (.Y(N9001),.A(N8501),.B(ttmp512));
OR2X1 OR2_2389 (.Y(N9005),.A(N4728),.B(N8516));
AND2X1 AND_tmp514 (.Y(ttmp514),.A(N6141),.B(N8537));
AND2X1 AND_tmp515 (.Y(N9024),.A(N7334),.B(ttmp514));
AND2X1 AND_tmp516 (.Y(ttmp516),.A(N7337),.B(N8538));
AND2X1 AND_tmp517 (.Y(N9025),.A(N6137),.B(ttmp516));
OR2X1 OR_tmp518 (.Y(ttmp518),.A(N8546),.B(N8547));
OR2X1 OR_tmp519 (.Y(ttmp519),.A(N4756),.B(ttmp518));
OR2X1 OR_tmp520 (.Y(N9029),.A(N8545),.B(ttmp519));
OR2X1 OR_tmp521 (.Y(ttmp521),.A(N8553),.B(N8554));
OR2X1 OR_tmp522 (.Y(ttmp522),.A(N4760),.B(ttmp521));
OR2X1 OR_tmp523 (.Y(ttmp523),.A(N8551),.B(ttmp522));
OR2X1 OR_tmp524 (.Y(N9035),.A(N8552),.B(ttmp523));
AND2X1 AND_tmp525 (.Y(ttmp525),.A(N6170),.B(N8564));
AND2X1 AND_tmp526 (.Y(N9053),.A(N7378),.B(ttmp525));
AND2X1 AND_tmp527 (.Y(ttmp527),.A(N7381),.B(N8565));
AND2X1 AND_tmp528 (.Y(N9054),.A(N6166),.B(ttmp527));
NAND2X1 NAND2_2396 (.Y(N9064),.A(N4303),.B(N8607));
NAND2X1 NAND2_2397 (.Y(N9065),.A(N3507),.B(N8609));
INVX1 NOT1_2398 (.Y(N9066),.A(N8114));
NAND2X1 NAND2_2399 (.Y(N9067),.A(N8114),.B(N4795));
OR2X1 OR2_2400 (.Y(N9068),.A(N7613),.B(N6783));
INVX1 NOT1_2401 (.Y(N9071),.A(N8117));
INVX1 NOT1_2402 (.Y(N9072),.A(N8131));
NAND2X1 NAND2_2403 (.Y(N9073),.A(N8131),.B(N6195));
INVX1 NOT1_2404 (.Y(N9074),.A(N7613));
INVX1 NOT1_2405 (.Y(N9077),.A(N8134));
OR2X1 OR2_2406 (.Y(N9079),.A(N7650),.B(N6865));
INVX1 NOT1_2407 (.Y(N9082),.A(N8146));
INVX1 NOT1_2408 (.Y(N9083),.A(N7650));
INVX1 NOT1_2409 (.Y(N9086),.A(N8156));
INVX1 NOT1_2410 (.Y(N9087),.A(N8166));
NAND2X1 NAND2_2411 (.Y(N9088),.A(N8166),.B(N4813));
OR2X1 OR2_2412 (.Y(N9089),.A(N7659),.B(N6866));
INVX1 NOT1_2413 (.Y(N9092),.A(N8169));
INVX1 NOT1_2414 (.Y(N9093),.A(N8183));
NAND2X1 NAND2_2415 (.Y(N9094),.A(N8183),.B(N6203));
INVX1 NOT1_2416 (.Y(N9095),.A(N7659));
INVX1 NOT1_2417 (.Y(N9098),.A(N8186));
OR2X1 OR_tmp529 (.Y(ttmp529),.A(N8341),.B(N8342));
OR2X1 OR_tmp530 (.Y(ttmp530),.A(N4545),.B(ttmp529));
OR2X1 OR_tmp531 (.Y(N9099),.A(N8340),.B(ttmp530));
OR2X1 OR_tmp532 (.Y(ttmp532),.A(N8343),.B(N8344));
NOR2X1 NOR_tmp533 (.Y(N9103),.A(N4545),.B(ttmp532));
OR2X1 OR_tmp534 (.Y(ttmp534),.A(N8345),.B(N8346));
OR2X1 OR_tmp535 (.Y(N9107),.A(N4549),.B(ttmp534));
NOR2X1 NOR2_2421 (.Y(N9111),.A(N4549),.B(N8347));
OR2X1 OR_tmp536 (.Y(ttmp536),.A(N8373),.B(N8374));
OR2X1 OR_tmp537 (.Y(ttmp537),.A(N4577),.B(ttmp536));
OR2X1 OR_tmp538 (.Y(N9117),.A(N8372),.B(ttmp537));
OR2X1 OR_tmp539 (.Y(ttmp539),.A(N8375),.B(N8376));
NOR2X1 NOR_tmp540 (.Y(N9127),.A(N4577),.B(ttmp539));
OR2X1 OR_tmp541 (.Y(ttmp541),.A(N8390),.B(N8391));
NOR2X1 NOR_tmp542 (.Y(N9146),.A(N4597),.B(ttmp541));
OR2X1 OR_tmp543 (.Y(ttmp543),.A(N8386),.B(N8387));
OR2X1 OR_tmp544 (.Y(ttmp544),.A(N4593),.B(ttmp543));
NOR2X1 NOR_tmp545 (.Y(N9149),.A(N8385),.B(ttmp544));
NAND2X1 NAND2_2426 (.Y(N9159),.A(N7577),.B(N8733));
NAND2X1 NAND2_2427 (.Y(N9160),.A(N7574),.B(N8734));
OR2X1 OR_tmp546 (.Y(ttmp546),.A(N8437),.B(N8438));
OR2X1 OR_tmp547 (.Y(ttmp547),.A(N4657),.B(ttmp546));
OR2X1 OR_tmp548 (.Y(N9161),.A(N8436),.B(ttmp547));
OR2X1 OR_tmp549 (.Y(ttmp549),.A(N8439),.B(N8440));
NOR2X1 NOR_tmp550 (.Y(N9165),.A(N4657),.B(ttmp549));
OR2X1 OR_tmp551 (.Y(ttmp551),.A(N8441),.B(N8442));
OR2X1 OR_tmp552 (.Y(N9169),.A(N4661),.B(ttmp551));
NOR2X1 NOR2_2431 (.Y(N9173),.A(N4661),.B(N8443));
NAND2X1 NAND2_2432 (.Y(N9179),.A(N7563),.B(N8753));
NAND2X1 NAND2_2433 (.Y(N9180),.A(N7560),.B(N8754));
NAND2X1 NAND2_2434 (.Y(N9181),.A(N7569),.B(N8755));
NAND2X1 NAND2_2435 (.Y(N9182),.A(N7566),.B(N8756));
OR2X1 OR_tmp553 (.Y(ttmp553),.A(N8492),.B(N8493));
OR2X1 OR_tmp554 (.Y(ttmp554),.A(N4702),.B(ttmp553));
OR2X1 OR_tmp555 (.Y(N9183),.A(N8491),.B(ttmp554));
OR2X1 OR_tmp556 (.Y(ttmp556),.A(N8494),.B(N8495));
NOR2X1 NOR_tmp557 (.Y(N9193),.A(N4702),.B(ttmp556));
OR2X1 OR_tmp558 (.Y(ttmp558),.A(N8512),.B(N8513));
OR2X1 OR_tmp559 (.Y(ttmp559),.A(N4722),.B(ttmp558));
OR2X1 OR_tmp560 (.Y(N9203),.A(N8511),.B(ttmp559));
OR2X1 OR_tmp561 (.Y(ttmp561),.A(N8506),.B(N8507));
OR2X1 OR_tmp562 (.Y(ttmp562),.A(N4718),.B(ttmp561));
OR2X1 OR_tmp563 (.Y(ttmp563),.A(N8504),.B(ttmp562));
OR2X1 OR_tmp564 (.Y(N9206),.A(N8505),.B(ttmp563));
OR2X1 OR_tmp565 (.Y(ttmp565),.A(N8514),.B(N8515));
NOR2X1 NOR_tmp566 (.Y(N9220),.A(N4722),.B(ttmp565));
OR2X1 OR_tmp567 (.Y(ttmp567),.A(N8509),.B(N8510));
OR2X1 OR_tmp568 (.Y(ttmp568),.A(N4718),.B(ttmp567));
NOR2X1 NOR_tmp569 (.Y(N9223),.A(N8508),.B(ttmp568));
NAND2X1 NAND2_2442 (.Y(N9234),.A(N7591),.B(N8814));
NAND2X1 NAND2_2443 (.Y(N9235),.A(N7588),.B(N8815));
NAND2X1 NAND2_2444 (.Y(N9236),.A(N7585),.B(N8816));
NAND2X1 NAND2_2445 (.Y(N9237),.A(N7582),.B(N8817));
OR2X1 OR2_2446 (.Y(N9238),.A(N3159),.B(N8818));
OR2X1 OR2_2447 (.Y(N9242),.A(N3126),.B(N8840));
NAND2X1 NAND2_2448 (.Y(N9243),.A(N8324),.B(N8888));
INVX1 NOT1_2449 (.Y(N9244),.A(N8580));
INVX1 NOT1_2450 (.Y(N9245),.A(N8583));
INVX1 NOT1_2451 (.Y(N9246),.A(N8586));
INVX1 NOT1_2452 (.Y(N9247),.A(N8589));
INVX1 NOT1_2453 (.Y(N9248),.A(N8592));
INVX1 NOT1_2454 (.Y(N9249),.A(N8595));
INVX1 NOT1_2455 (.Y(N9250),.A(N8598));
INVX1 NOT1_2456 (.Y(N9251),.A(N8601));
INVX1 NOT1_2457 (.Y(N9252),.A(N8604));
NOR2X1 NOR2_2458 (.Y(N9256),.A(N8861),.B(N8280));
NOR2X1 NOR2_2459 (.Y(N9257),.A(N8862),.B(N8281));
NOR2X1 NOR2_2460 (.Y(N9258),.A(N8863),.B(N8282));
NOR2X1 NOR2_2461 (.Y(N9259),.A(N8864),.B(N8283));
NOR2X1 NOR2_2462 (.Y(N9260),.A(N8865),.B(N8284));
NOR2X1 NOR2_2463 (.Y(N9261),.A(N8866),.B(N8285));
INVX1 NOT1_2464 (.Y(N9262),.A(N8627));
OR2X1 OR2_2465 (.Y(N9265),.A(N7649),.B(N8874));
OR2X1 OR2_2466 (.Y(N9268),.A(N7668),.B(N8878));
NAND2X1 NAND2_2467 (.Y(N9271),.A(N7533),.B(N8879));
NAND2X1 NAND2_2468 (.Y(N9272),.A(N7536),.B(N8881));
NAND2X1 NAND2_2469 (.Y(N9273),.A(N7539),.B(N8883));
NAND2X1 NAND2_2470 (.Y(N9274),.A(N7542),.B(N8885));
NAND2X1 NAND2_2471 (.Y(N9275),.A(N8322),.B(N8887));
INVX1 NOT1_2472 (.Y(N9276),.A(N8333));
AND2X1 AND_tmp570 (.Y(ttmp570),.A(N6929),.B(N6957));
AND2X1 AND_tmp571 (.Y(ttmp571),.A(N6936),.B(ttmp570));
AND2X1 AND_tmp572 (.Y(ttmp572),.A(N8326),.B(ttmp571));
AND2X1 AND_tmp573 (.Y(N9280),.A(N6946),.B(ttmp572));
AND2X1 AND_tmp574 (.Y(ttmp574),.A(N6957),.B(N6936));
AND2X1 AND_tmp575 (.Y(ttmp575),.A(N367),.B(ttmp574));
AND2X1 AND_tmp576 (.Y(ttmp576),.A(N8326),.B(ttmp575));
AND2X1 AND_tmp577 (.Y(N9285),.A(N6946),.B(ttmp576));
AND2X1 AND_tmp578 (.Y(ttmp578),.A(N6946),.B(N6957));
AND2X1 AND_tmp579 (.Y(ttmp579),.A(N367),.B(ttmp578));
AND2X1 AND_tmp580 (.Y(N9286),.A(N8326),.B(ttmp579));
AND2X1 AND_tmp581 (.Y(ttmp581),.A(N8326),.B(N6957));
AND2X1 AND_tmp582 (.Y(N9287),.A(N367),.B(ttmp581));
AND2X1 AND2_2477 (.Y(N9288),.A(N367),.B(N8326));
INVX1 NOT1_2478 (.Y(N9290),.A(N8660));
INVX1 NOT1_2479 (.Y(N9292),.A(N8663));
INVX1 NOT1_2480 (.Y(N9294),.A(N8666));
INVX1 NOT1_2481 (.Y(N9296),.A(N8669));
NAND2X1 NAND2_2482 (.Y(N9297),.A(N8672),.B(N5966));
INVX1 NOT1_2483 (.Y(N9298),.A(N8672));
NAND2X1 NAND2_2484 (.Y(N9299),.A(N8675),.B(N6969));
INVX1 NOT1_2485 (.Y(N9300),.A(N8675));
INVX1 NOT1_2486 (.Y(N9301),.A(N8365));
AND2X1 AND_tmp583 (.Y(ttmp583),.A(N7006),.B(N6998));
AND2X1 AND_tmp584 (.Y(ttmp584),.A(N8358),.B(ttmp583));
AND2X1 AND_tmp585 (.Y(ttmp585),.A(N7036),.B(ttmp584));
AND2X1 AND_tmp586 (.Y(N9307),.A(N7020),.B(ttmp585));
AND2X1 AND_tmp587 (.Y(ttmp587),.A(N7006),.B(N7036));
AND2X1 AND_tmp588 (.Y(ttmp588),.A(N8358),.B(ttmp587));
AND2X1 AND_tmp589 (.Y(N9314),.A(N7020),.B(ttmp588));
AND2X1 AND_tmp590 (.Y(ttmp590),.A(N7020),.B(N7036));
AND2X1 AND_tmp591 (.Y(N9315),.A(N8358),.B(ttmp590));
AND2X1 AND2_2490 (.Y(N9318),.A(N8358),.B(N7036));
INVX1 NOT1_2491 (.Y(N9319),.A(N8687));
INVX1 NOT1_2492 (.Y(N9320),.A(N8699));
INVX1 NOT1_2493 (.Y(N9321),.A(N8711));
INVX1 NOT1_2494 (.Y(N9322),.A(N8714));
INVX1 NOT1_2495 (.Y(N9323),.A(N8727));
INVX1 NOT1_2496 (.Y(N9324),.A(N8730));
INVX1 NOT1_2497 (.Y(N9326),.A(N8405));
AND2X1 AND2_2498 (.Y(N9332),.A(N8405),.B(N8412));
OR2X1 OR2_2499 (.Y(N9339),.A(N4193),.B(N8960));
AND2X1 AND2_2500 (.Y(N9344),.A(N8430),.B(N8444));
INVX1 NOT1_2501 (.Y(N9352),.A(N8735));
INVX1 NOT1_2502 (.Y(N9354),.A(N8738));
INVX1 NOT1_2503 (.Y(N9356),.A(N8741));
INVX1 NOT1_2504 (.Y(N9358),.A(N8744));
NAND2X1 NAND2_2505 (.Y(N9359),.A(N8747),.B(N6078));
INVX1 NOT1_2506 (.Y(N9360),.A(N8747));
NAND2X1 NAND2_2507 (.Y(N9361),.A(N8750),.B(N7187));
INVX1 NOT1_2508 (.Y(N9362),.A(N8750));
INVX1 NOT1_2509 (.Y(N9363),.A(N8471));
INVX1 NOT1_2510 (.Y(N9364),.A(N8474));
INVX1 NOT1_2511 (.Y(N9365),.A(N8477));
INVX1 NOT1_2512 (.Y(N9366),.A(N8480));
NOR2X1 NOR2_2513 (.Y(N9367),.A(N8991),.B(N8483));
NOR2X1 NOR2_2514 (.Y(N9368),.A(N8992),.B(N8484));
AND2X1 AND_tmp592 (.Y(ttmp592),.A(N7194),.B(N8471));
AND2X1 AND_tmp593 (.Y(N9369),.A(N7198),.B(ttmp592));
AND2X1 AND_tmp594 (.Y(ttmp594),.A(N8457),.B(N8474));
AND2X1 AND_tmp595 (.Y(N9370),.A(N8460),.B(ttmp594));
AND2X1 AND_tmp596 (.Y(ttmp596),.A(N7205),.B(N8477));
AND2X1 AND_tmp597 (.Y(N9371),.A(N7209),.B(ttmp596));
AND2X1 AND_tmp598 (.Y(ttmp598),.A(N8463),.B(N8480));
AND2X1 AND_tmp599 (.Y(N9372),.A(N8466),.B(ttmp598));
INVX1 NOT1_2519 (.Y(N9375),.A(N8497));
INVX1 NOT1_2520 (.Y(N9381),.A(N8766));
INVX1 NOT1_2521 (.Y(N9382),.A(N8778));
INVX1 NOT1_2522 (.Y(N9383),.A(N8793));
INVX1 NOT1_2523 (.Y(N9384),.A(N8796));
AND2X1 AND2_2524 (.Y(N9385),.A(N8485),.B(N8497));
INVX1 NOT1_2525 (.Y(N9392),.A(N8525));
INVX1 NOT1_2526 (.Y(N9393),.A(N8528));
INVX1 NOT1_2527 (.Y(N9394),.A(N8531));
INVX1 NOT1_2528 (.Y(N9395),.A(N8534));
AND2X1 AND_tmp600 (.Y(ttmp600),.A(N7314),.B(N8525));
AND2X1 AND_tmp601 (.Y(N9396),.A(N7318),.B(ttmp600));
AND2X1 AND_tmp602 (.Y(ttmp602),.A(N8519),.B(N8528));
AND2X1 AND_tmp603 (.Y(N9397),.A(N8522),.B(ttmp602));
AND2X1 AND_tmp604 (.Y(ttmp604),.A(N6127),.B(N8531));
AND2X1 AND_tmp605 (.Y(N9398),.A(N6131),.B(ttmp604));
AND2X1 AND_tmp606 (.Y(ttmp606),.A(N7325),.B(N8534));
AND2X1 AND_tmp607 (.Y(N9399),.A(N7328),.B(ttmp606));
NOR2X1 NOR2_2533 (.Y(N9400),.A(N9024),.B(N8539));
NOR2X1 NOR2_2534 (.Y(N9401),.A(N9025),.B(N8540));
INVX1 NOT1_2535 (.Y(N9402),.A(N8541));
NAND2X1 NAND2_2536 (.Y(N9407),.A(N8548),.B(N89));
AND2X1 AND2_2537 (.Y(N9408),.A(N8541),.B(N8548));
INVX1 NOT1_2538 (.Y(N9412),.A(N8811));
INVX1 NOT1_2539 (.Y(N9413),.A(N8566));
INVX1 NOT1_2540 (.Y(N9414),.A(N8569));
INVX1 NOT1_2541 (.Y(N9415),.A(N8572));
INVX1 NOT1_2542 (.Y(N9416),.A(N8575));
NOR2X1 NOR2_2543 (.Y(N9417),.A(N9053),.B(N8578));
NOR2X1 NOR2_2544 (.Y(N9418),.A(N9054),.B(N8579));
AND2X1 AND_tmp608 (.Y(ttmp608),.A(N6177),.B(N8566));
AND2X1 AND_tmp609 (.Y(N9419),.A(N7387),.B(ttmp608));
AND2X1 AND_tmp610 (.Y(ttmp610),.A(N7384),.B(N8569));
AND2X1 AND_tmp611 (.Y(N9420),.A(N8555),.B(ttmp610));
AND2X1 AND_tmp612 (.Y(ttmp612),.A(N7394),.B(N8572));
AND2X1 AND_tmp613 (.Y(N9421),.A(N7398),.B(ttmp612));
AND2X1 AND_tmp614 (.Y(ttmp614),.A(N8558),.B(N8575));
AND2X1 AND_tmp615 (.Y(N9422),.A(N8561),.B(ttmp614));
BUFX1 BUFF1_2549 (.Y(N9423),.A(N8326));
NAND2X1 NAND2_2550 (.Y(N9426),.A(N9064),.B(N8608));
NAND2X1 NAND2_2551 (.Y(N9429),.A(N9065),.B(N8610));
NAND2X1 NAND2_2552 (.Y(N9432),.A(N3515),.B(N9066));
NAND2X1 NAND2_2553 (.Y(N9435),.A(N4796),.B(N9072));
NAND2X1 NAND2_2554 (.Y(N9442),.A(N3628),.B(N9087));
NAND2X1 NAND2_2555 (.Y(N9445),.A(N4814),.B(N9093));
INVX1 NOT1_2556 (.Y(N9454),.A(N8678));
INVX1 NOT1_2557 (.Y(N9455),.A(N8681));
INVX1 NOT1_2558 (.Y(N9456),.A(N8684));
INVX1 NOT1_2559 (.Y(N9459),.A(N8690));
INVX1 NOT1_2560 (.Y(N9460),.A(N8693));
INVX1 NOT1_2561 (.Y(N9461),.A(N8696));
BUFX1 BUFF1_2562 (.Y(N9462),.A(N8358));
INVX1 NOT1_2563 (.Y(N9465),.A(N8702));
INVX1 NOT1_2564 (.Y(N9466),.A(N8705));
INVX1 NOT1_2565 (.Y(N9467),.A(N8708));
INVX1 NOT1_2566 (.Y(N9468),.A(N8724));
BUFX1 BUFF1_2567 (.Y(N9473),.A(N8358));
INVX1 NOT1_2568 (.Y(N9476),.A(N8718));
INVX1 NOT1_2569 (.Y(N9477),.A(N8721));
NAND2X1 NAND2_2570 (.Y(N9478),.A(N9159),.B(N9160));
NAND2X1 NAND2_2571 (.Y(N9485),.A(N9179),.B(N9180));
NAND2X1 NAND2_2572 (.Y(N9488),.A(N9181),.B(N9182));
INVX1 NOT1_2573 (.Y(N9493),.A(N8757));
INVX1 NOT1_2574 (.Y(N9494),.A(N8760));
INVX1 NOT1_2575 (.Y(N9495),.A(N8763));
INVX1 NOT1_2576 (.Y(N9498),.A(N8769));
INVX1 NOT1_2577 (.Y(N9499),.A(N8772));
INVX1 NOT1_2578 (.Y(N9500),.A(N8775));
INVX1 NOT1_2579 (.Y(N9505),.A(N8781));
INVX1 NOT1_2580 (.Y(N9506),.A(N8784));
INVX1 NOT1_2581 (.Y(N9507),.A(N8787));
INVX1 NOT1_2582 (.Y(N9508),.A(N8790));
INVX1 NOT1_2583 (.Y(N9509),.A(N8808));
INVX1 NOT1_2584 (.Y(N9514),.A(N8799));
INVX1 NOT1_2585 (.Y(N9515),.A(N8802));
INVX1 NOT1_2586 (.Y(N9516),.A(N8805));
NAND2X1 NAND2_2587 (.Y(N9517),.A(N9234),.B(N9235));
NAND2X1 NAND2_2588 (.Y(N9520),.A(N9236),.B(N9237));
AND2X1 AND2_2589 (.Y(N9526),.A(N8943),.B(N8421));
AND2X1 AND2_2590 (.Y(N9531),.A(N8943),.B(N8421));
NAND2X1 NAND2_2591 (.Y(N9539),.A(N9271),.B(N8880));
NAND2X1 NAND2_2592 (.Y(N9540),.A(N9273),.B(N8884));
INVX1 NOT1_2593 (.Y(N9541),.A(N9275));
AND2X1 AND2_2594 (.Y(N9543),.A(N8857),.B(N8254));
AND2X1 AND2_2595 (.Y(N9551),.A(N8871),.B(N8288));
NAND2X1 NAND2_2596 (.Y(N9555),.A(N9272),.B(N8882));
NAND2X1 NAND2_2597 (.Y(N9556),.A(N9274),.B(N8886));
INVX1 NOT1_2598 (.Y(N9557),.A(N8898));
AND2X1 AND2_2599 (.Y(N9560),.A(N8902),.B(N8333));
INVX1 NOT1_2600 (.Y(N9561),.A(N9099));
NAND2X1 NAND2_2601 (.Y(N9562),.A(N9099),.B(N9290));
INVX1 NOT1_2602 (.Y(N9563),.A(N9103));
NAND2X1 NAND2_2603 (.Y(N9564),.A(N9103),.B(N9292));
INVX1 NOT1_2604 (.Y(N9565),.A(N9107));
NAND2X1 NAND2_2605 (.Y(N9566),.A(N9107),.B(N9294));
INVX1 NOT1_2606 (.Y(N9567),.A(N9111));
NAND2X1 NAND2_2607 (.Y(N9568),.A(N9111),.B(N9296));
NAND2X1 NAND2_2608 (.Y(N9569),.A(N4844),.B(N9298));
NAND2X1 NAND2_2609 (.Y(N9570),.A(N6207),.B(N9300));
INVX1 NOT1_2610 (.Y(N9571),.A(N8920));
INVX1 NOT1_2611 (.Y(N9575),.A(N8927));
AND2X1 AND2_2612 (.Y(N9579),.A(N8365),.B(N8927));
INVX1 NOT1_2613 (.Y(N9581),.A(N8950));
INVX1 NOT1_2614 (.Y(N9582),.A(N8956));
AND2X1 AND2_2615 (.Y(N9585),.A(N8405),.B(N8956));
AND2X1 AND2_2616 (.Y(N9591),.A(N8966),.B(N8430));
INVX1 NOT1_2617 (.Y(N9592),.A(N9161));
NAND2X1 NAND2_2618 (.Y(N9593),.A(N9161),.B(N9352));
INVX1 NOT1_2619 (.Y(N9594),.A(N9165));
NAND2X1 NAND2_2620 (.Y(N9595),.A(N9165),.B(N9354));
INVX1 NOT1_2621 (.Y(N9596),.A(N9169));
NAND2X1 NAND2_2622 (.Y(N9597),.A(N9169),.B(N9356));
INVX1 NOT1_2623 (.Y(N9598),.A(N9173));
NAND2X1 NAND2_2624 (.Y(N9599),.A(N9173),.B(N9358));
NAND2X1 NAND2_2625 (.Y(N9600),.A(N4940),.B(N9360));
NAND2X1 NAND2_2626 (.Y(N9601),.A(N6220),.B(N9362));
AND2X1 AND_tmp616 (.Y(ttmp616),.A(N7198),.B(N9363));
AND2X1 AND_tmp617 (.Y(N9602),.A(N8457),.B(ttmp616));
AND2X1 AND_tmp618 (.Y(ttmp618),.A(N8460),.B(N9364));
AND2X1 AND_tmp619 (.Y(N9603),.A(N7194),.B(ttmp618));
AND2X1 AND_tmp620 (.Y(ttmp620),.A(N7209),.B(N9365));
AND2X1 AND_tmp621 (.Y(N9604),.A(N8463),.B(ttmp620));
AND2X1 AND_tmp622 (.Y(ttmp622),.A(N8466),.B(N9366));
AND2X1 AND_tmp623 (.Y(N9605),.A(N7205),.B(ttmp622));
INVX1 NOT1_2631 (.Y(N9608),.A(N9001));
AND2X1 AND2_2632 (.Y(N9611),.A(N8485),.B(N9001));
AND2X1 AND_tmp624 (.Y(ttmp624),.A(N7318),.B(N9392));
AND2X1 AND_tmp625 (.Y(N9612),.A(N8519),.B(ttmp624));
AND2X1 AND_tmp626 (.Y(ttmp626),.A(N8522),.B(N9393));
AND2X1 AND_tmp627 (.Y(N9613),.A(N7314),.B(ttmp626));
AND2X1 AND_tmp628 (.Y(ttmp628),.A(N6131),.B(N9394));
AND2X1 AND_tmp629 (.Y(N9614),.A(N7325),.B(ttmp628));
AND2X1 AND_tmp630 (.Y(ttmp630),.A(N7328),.B(N9395));
AND2X1 AND_tmp631 (.Y(N9615),.A(N6127),.B(ttmp630));
INVX1 NOT1_2637 (.Y(N9616),.A(N9029));
INVX1 NOT1_2638 (.Y(N9617),.A(N9035));
AND2X1 AND2_2639 (.Y(N9618),.A(N8541),.B(N9035));
AND2X1 AND_tmp632 (.Y(ttmp632),.A(N7387),.B(N9413));
AND2X1 AND_tmp633 (.Y(N9621),.A(N7384),.B(ttmp632));
AND2X1 AND_tmp634 (.Y(ttmp634),.A(N8555),.B(N9414));
AND2X1 AND_tmp635 (.Y(N9622),.A(N6177),.B(ttmp634));
AND2X1 AND_tmp636 (.Y(ttmp636),.A(N7398),.B(N9415));
AND2X1 AND_tmp637 (.Y(N9623),.A(N8558),.B(ttmp636));
AND2X1 AND_tmp638 (.Y(ttmp638),.A(N8561),.B(N9416));
AND2X1 AND_tmp639 (.Y(N9624),.A(N7394),.B(ttmp638));
OR2X1 OR_tmp640 (.Y(ttmp640),.A(N8354),.B(N9285));
OR2X1 OR_tmp641 (.Y(ttmp641),.A(N4563),.B(ttmp640));
OR2X1 OR_tmp642 (.Y(ttmp642),.A(N8352),.B(ttmp641));
OR2X1 OR_tmp643 (.Y(N9626),.A(N8353),.B(ttmp642));
OR2X1 OR_tmp644 (.Y(ttmp644),.A(N8356),.B(N9286));
OR2X1 OR_tmp645 (.Y(ttmp645),.A(N4566),.B(ttmp644));
OR2X1 OR_tmp646 (.Y(N9629),.A(N8355),.B(ttmp645));
OR2X1 OR_tmp647 (.Y(ttmp647),.A(N8357),.B(N9287));
OR2X1 OR_tmp648 (.Y(N9632),.A(N4570),.B(ttmp647));
OR2X1 OR2_2647 (.Y(N9635),.A(N5960),.B(N9288));
NAND2X1 NAND2_2648 (.Y(N9642),.A(N9067),.B(N9432));
INVX1 NOT1_2649 (.Y(N9645),.A(N9068));
NAND2X1 NAND2_2650 (.Y(N9646),.A(N9073),.B(N9435));
INVX1 NOT1_2651 (.Y(N9649),.A(N9074));
NAND2X1 NAND2_2652 (.Y(N9650),.A(N9257),.B(N9256));
NAND2X1 NAND2_2653 (.Y(N9653),.A(N9259),.B(N9258));
NAND2X1 NAND2_2654 (.Y(N9656),.A(N9261),.B(N9260));
INVX1 NOT1_2655 (.Y(N9659),.A(N9079));
NAND2X1 NAND2_2656 (.Y(N9660),.A(N9079),.B(N4809));
INVX1 NOT1_2657 (.Y(N9661),.A(N9083));
NAND2X1 NAND2_2658 (.Y(N9662),.A(N9083),.B(N6202));
NAND2X1 NAND2_2659 (.Y(N9663),.A(N9088),.B(N9442));
INVX1 NOT1_2660 (.Y(N9666),.A(N9089));
NAND2X1 NAND2_2661 (.Y(N9667),.A(N9094),.B(N9445));
INVX1 NOT1_2662 (.Y(N9670),.A(N9095));
OR2X1 OR2_2663 (.Y(N9671),.A(N8924),.B(N8393));
INVX1 NOT1_2664 (.Y(N9674),.A(N9117));
INVX1 NOT1_2665 (.Y(N9675),.A(N8924));
INVX1 NOT1_2666 (.Y(N9678),.A(N9127));
OR2X1 OR_tmp649 (.Y(ttmp649),.A(N8389),.B(N9315));
OR2X1 OR_tmp650 (.Y(ttmp650),.A(N4597),.B(ttmp649));
OR2X1 OR_tmp651 (.Y(N9679),.A(N8388),.B(ttmp650));
OR2X1 OR2_2668 (.Y(N9682),.A(N8931),.B(N9318));
OR2X1 OR_tmp652 (.Y(ttmp652),.A(N8384),.B(N9314));
OR2X1 OR_tmp653 (.Y(ttmp653),.A(N4593),.B(ttmp652));
OR2X1 OR_tmp654 (.Y(ttmp654),.A(N8382),.B(ttmp653));
OR2X1 OR_tmp655 (.Y(N9685),.A(N8383),.B(ttmp654));
INVX1 NOT1_2670 (.Y(N9690),.A(N9146));
NAND2X1 NAND2_2671 (.Y(N9691),.A(N9146),.B(N8717));
INVX1 NOT1_2672 (.Y(N9692),.A(N8931));
INVX1 NOT1_2673 (.Y(N9695),.A(N9149));
NAND2X1 NAND2_2674 (.Y(N9698),.A(N9401),.B(N9400));
NAND2X1 NAND2_2675 (.Y(N9702),.A(N9368),.B(N9367));
OR2X1 OR2_2676 (.Y(N9707),.A(N8996),.B(N8517));
INVX1 NOT1_2677 (.Y(N9710),.A(N9183));
INVX1 NOT1_2678 (.Y(N9711),.A(N8996));
INVX1 NOT1_2679 (.Y(N9714),.A(N9193));
INVX1 NOT1_2680 (.Y(N9715),.A(N9203));
NAND2X1 NAND2_2681 (.Y(N9716),.A(N9203),.B(N6235));
OR2X1 OR2_2682 (.Y(N9717),.A(N9005),.B(N8518));
INVX1 NOT1_2683 (.Y(N9720),.A(N9206));
INVX1 NOT1_2684 (.Y(N9721),.A(N9220));
NAND2X1 NAND2_2685 (.Y(N9722),.A(N9220),.B(N7573));
INVX1 NOT1_2686 (.Y(N9723),.A(N9005));
INVX1 NOT1_2687 (.Y(N9726),.A(N9223));
NAND2X1 NAND2_2688 (.Y(N9727),.A(N9418),.B(N9417));
AND2X1 AND2_2689 (.Y(N9732),.A(N9268),.B(N8269));
NAND2X1 NAND2_2690 (.Y(N9733),.A(N9581),.B(N9326));
AND2X1 AND_tmp656 (.Y(ttmp656),.A(N8394),.B(N8421));
AND2X1 AND_tmp657 (.Y(ttmp657),.A(N89),.B(ttmp656));
AND2X1 AND_tmp658 (.Y(ttmp658),.A(N9408),.B(ttmp657));
AND2X1 AND_tmp659 (.Y(N9734),.A(N9332),.B(ttmp658));
AND2X1 AND_tmp660 (.Y(ttmp660),.A(N8394),.B(N8421));
AND2X1 AND_tmp661 (.Y(ttmp661),.A(N89),.B(ttmp660));
AND2X1 AND_tmp662 (.Y(ttmp662),.A(N9408),.B(ttmp661));
AND2X1 AND_tmp663 (.Y(N9735),.A(N9332),.B(ttmp662));
AND2X1 AND2_2693 (.Y(N9736),.A(N9265),.B(N8262));
INVX1 NOT1_2694 (.Y(N9737),.A(N9555));
INVX1 NOT1_2695 (.Y(N9738),.A(N9556));
NAND2X1 NAND2_2696 (.Y(N9739),.A(N9361),.B(N9601));
NAND2X1 NAND2_2697 (.Y(N9740),.A(N9423),.B(N1115));
INVX1 NOT1_2698 (.Y(N9741),.A(N9423));
NAND2X1 NAND2_2699 (.Y(N9742),.A(N9299),.B(N9570));
AND2X1 AND2_2700 (.Y(N9754),.A(N8333),.B(N9280));
OR2X1 OR2_2701 (.Y(N9758),.A(N8898),.B(N9560));
NAND2X1 NAND2_2702 (.Y(N9762),.A(N8660),.B(N9561));
NAND2X1 NAND2_2703 (.Y(N9763),.A(N8663),.B(N9563));
NAND2X1 NAND2_2704 (.Y(N9764),.A(N8666),.B(N9565));
NAND2X1 NAND2_2705 (.Y(N9765),.A(N8669),.B(N9567));
NAND2X1 NAND2_2706 (.Y(N9766),.A(N9297),.B(N9569));
AND2X1 AND2_2707 (.Y(N9767),.A(N9280),.B(N367));
NAND2X1 NAND2_2708 (.Y(N9768),.A(N9557),.B(N9276));
INVX1 NOT1_2709 (.Y(N9769),.A(N9307));
NAND2X1 NAND2_2710 (.Y(N9773),.A(N9307),.B(N367));
NAND2X1 NAND2_2711 (.Y(N9774),.A(N9571),.B(N9301));
AND2X1 AND2_2712 (.Y(N9775),.A(N8365),.B(N9307));
OR2X1 OR2_2713 (.Y(N9779),.A(N8920),.B(N9579));
INVX1 NOT1_2714 (.Y(N9784),.A(N9478));
NAND2X1 NAND2_2715 (.Y(N9785),.A(N9616),.B(N9402));
OR2X1 OR2_2716 (.Y(N9786),.A(N8950),.B(N9585));
AND2X1 AND_tmp664 (.Y(ttmp664),.A(N9332),.B(N8394));
AND2X1 AND_tmp665 (.Y(ttmp665),.A(N89),.B(ttmp664));
AND2X1 AND_tmp666 (.Y(N9790),.A(N9408),.B(ttmp665));
OR2X1 OR2_2718 (.Y(N9791),.A(N8963),.B(N9591));
NAND2X1 NAND2_2719 (.Y(N9795),.A(N8735),.B(N9592));
NAND2X1 NAND2_2720 (.Y(N9796),.A(N8738),.B(N9594));
NAND2X1 NAND2_2721 (.Y(N9797),.A(N8741),.B(N9596));
NAND2X1 NAND2_2722 (.Y(N9798),.A(N8744),.B(N9598));
NAND2X1 NAND2_2723 (.Y(N9799),.A(N9359),.B(N9600));
NOR2X1 NOR2_2724 (.Y(N9800),.A(N9602),.B(N9369));
NOR2X1 NOR2_2725 (.Y(N9801),.A(N9603),.B(N9370));
NOR2X1 NOR2_2726 (.Y(N9802),.A(N9604),.B(N9371));
NOR2X1 NOR2_2727 (.Y(N9803),.A(N9605),.B(N9372));
INVX1 NOT1_2728 (.Y(N9805),.A(N9485));
INVX1 NOT1_2729 (.Y(N9806),.A(N9488));
OR2X1 OR2_2730 (.Y(N9809),.A(N8995),.B(N9611));
NOR2X1 NOR2_2731 (.Y(N9813),.A(N9612),.B(N9396));
NOR2X1 NOR2_2732 (.Y(N9814),.A(N9613),.B(N9397));
NOR2X1 NOR2_2733 (.Y(N9815),.A(N9614),.B(N9398));
NOR2X1 NOR2_2734 (.Y(N9816),.A(N9615),.B(N9399));
AND2X1 AND2_2735 (.Y(N9817),.A(N9617),.B(N9407));
OR2X1 OR2_2736 (.Y(N9820),.A(N9029),.B(N9618));
INVX1 NOT1_2737 (.Y(N9825),.A(N9517));
INVX1 NOT1_2738 (.Y(N9826),.A(N9520));
NOR2X1 NOR2_2739 (.Y(N9827),.A(N9621),.B(N9419));
NOR2X1 NOR2_2740 (.Y(N9828),.A(N9622),.B(N9420));
NOR2X1 NOR2_2741 (.Y(N9829),.A(N9623),.B(N9421));
NOR2X1 NOR2_2742 (.Y(N9830),.A(N9624),.B(N9422));
INVX1 NOT1_2743 (.Y(N9835),.A(N9426));
NAND2X1 NAND2_2744 (.Y(N9836),.A(N9426),.B(N4789));
INVX1 NOT1_2745 (.Y(N9837),.A(N9429));
NAND2X1 NAND2_2746 (.Y(N9838),.A(N9429),.B(N4794));
NAND2X1 NAND2_2747 (.Y(N9846),.A(N3625),.B(N9659));
NAND2X1 NAND2_2748 (.Y(N9847),.A(N4810),.B(N9661));
INVX1 NOT1_2749 (.Y(N9862),.A(N9462));
NAND2X1 NAND2_2750 (.Y(N9863),.A(N7553),.B(N9690));
INVX1 NOT1_2751 (.Y(N9866),.A(N9473));
NAND2X1 NAND2_2752 (.Y(N9873),.A(N5030),.B(N9715));
NAND2X1 NAND2_2753 (.Y(N9876),.A(N6236),.B(N9721));
NAND2X1 NAND2_2754 (.Y(N9890),.A(N9795),.B(N9593));
NAND2X1 NAND2_2755 (.Y(N9891),.A(N9797),.B(N9597));
INVX1 NOT1_2756 (.Y(N9892),.A(N9799));
NAND2X1 NAND2_2757 (.Y(N9893),.A(N871),.B(N9741));
NAND2X1 NAND2_2758 (.Y(N9894),.A(N9762),.B(N9562));
NAND2X1 NAND2_2759 (.Y(N9895),.A(N9764),.B(N9566));
INVX1 NOT1_2760 (.Y(N9896),.A(N9766));
INVX1 NOT1_2761 (.Y(N9897),.A(N9626));
NAND2X1 NAND2_2762 (.Y(N9898),.A(N9626),.B(N9249));
INVX1 NOT1_2763 (.Y(N9899),.A(N9629));
NAND2X1 NAND2_2764 (.Y(N9900),.A(N9629),.B(N9250));
INVX1 NOT1_2765 (.Y(N9901),.A(N9632));
NAND2X1 NAND2_2766 (.Y(N9902),.A(N9632),.B(N9251));
INVX1 NOT1_2767 (.Y(N9903),.A(N9635));
NAND2X1 NAND2_2768 (.Y(N9904),.A(N9635),.B(N9252));
INVX1 NOT1_2769 (.Y(N9905),.A(N9543));
INVX1 NOT1_2770 (.Y(N9906),.A(N9650));
NAND2X1 NAND2_2771 (.Y(N9907),.A(N9650),.B(N5769));
INVX1 NOT1_2772 (.Y(N9908),.A(N9653));
NAND2X1 NAND2_2773 (.Y(N9909),.A(N9653),.B(N5770));
INVX1 NOT1_2774 (.Y(N9910),.A(N9656));
NAND2X1 NAND2_2775 (.Y(N9911),.A(N9656),.B(N9262));
INVX1 NOT1_2776 (.Y(N9917),.A(N9551));
NAND2X1 NAND2_2777 (.Y(N9923),.A(N9763),.B(N9564));
NAND2X1 NAND2_2778 (.Y(N9924),.A(N9765),.B(N9568));
OR2X1 OR2_2779 (.Y(N9925),.A(N8902),.B(N9767));
AND2X1 AND2_2780 (.Y(N9932),.A(N9575),.B(N9773));
AND2X1 AND2_2781 (.Y(N9935),.A(N9575),.B(N9769));
INVX1 NOT1_2782 (.Y(N9938),.A(N9698));
NAND2X1 NAND2_2783 (.Y(N9939),.A(N9698),.B(N9323));
NAND2X1 NAND2_2784 (.Y(N9945),.A(N9796),.B(N9595));
NAND2X1 NAND2_2785 (.Y(N9946),.A(N9798),.B(N9599));
INVX1 NOT1_2786 (.Y(N9947),.A(N9702));
NAND2X1 NAND2_2787 (.Y(N9948),.A(N9702),.B(N6102));
AND2X1 AND2_2788 (.Y(N9949),.A(N9608),.B(N9375));
INVX1 NOT1_2789 (.Y(N9953),.A(N9727));
NAND2X1 NAND2_2790 (.Y(N9954),.A(N9727),.B(N9412));
NAND2X1 NAND2_2791 (.Y(N9955),.A(N3502),.B(N9835));
NAND2X1 NAND2_2792 (.Y(N9956),.A(N3510),.B(N9837));
INVX1 NOT1_2793 (.Y(N9957),.A(N9642));
NAND2X1 NAND2_2794 (.Y(N9958),.A(N9642),.B(N9645));
INVX1 NOT1_2795 (.Y(N9959),.A(N9646));
NAND2X1 NAND2_2796 (.Y(N9960),.A(N9646),.B(N9649));
NAND2X1 NAND2_2797 (.Y(N9961),.A(N9660),.B(N9846));
NAND2X1 NAND2_2798 (.Y(N9964),.A(N9662),.B(N9847));
INVX1 NOT1_2799 (.Y(N9967),.A(N9663));
NAND2X1 NAND2_2800 (.Y(N9968),.A(N9663),.B(N9666));
INVX1 NOT1_2801 (.Y(N9969),.A(N9667));
NAND2X1 NAND2_2802 (.Y(N9970),.A(N9667),.B(N9670));
INVX1 NOT1_2803 (.Y(N9971),.A(N9671));
NAND2X1 NAND2_2804 (.Y(N9972),.A(N9671),.B(N6213));
INVX1 NOT1_2805 (.Y(N9973),.A(N9675));
NAND2X1 NAND2_2806 (.Y(N9974),.A(N9675),.B(N7551));
INVX1 NOT1_2807 (.Y(N9975),.A(N9679));
NAND2X1 NAND2_2808 (.Y(N9976),.A(N9679),.B(N7552));
INVX1 NOT1_2809 (.Y(N9977),.A(N9682));
INVX1 NOT1_2810 (.Y(N9978),.A(N9685));
NAND2X1 NAND2_2811 (.Y(N9979),.A(N9691),.B(N9863));
INVX1 NOT1_2812 (.Y(N9982),.A(N9692));
NAND2X1 NAND2_2813 (.Y(N9983),.A(N9814),.B(N9813));
NAND2X1 NAND2_2814 (.Y(N9986),.A(N9816),.B(N9815));
NAND2X1 NAND2_2815 (.Y(N9989),.A(N9801),.B(N9800));
NAND2X1 NAND2_2816 (.Y(N9992),.A(N9803),.B(N9802));
INVX1 NOT1_2817 (.Y(N9995),.A(N9707));
NAND2X1 NAND2_2818 (.Y(N9996),.A(N9707),.B(N6231));
INVX1 NOT1_2819 (.Y(N9997),.A(N9711));
NAND2X1 NAND2_2820 (.Y(N9998),.A(N9711),.B(N7572));
NAND2X1 NAND2_2821 (.Y(N9999),.A(N9716),.B(N9873));
INVX1 NOT1_2822 (.Y(N10002),.A(N9717));
NAND2X1 NAND2_2823 (.Y(N10003),.A(N9722),.B(N9876));
INVX1 NOT1_2824 (.Y(N10006),.A(N9723));
NAND2X1 NAND2_2825 (.Y(N10007),.A(N9830),.B(N9829));
NAND2X1 NAND2_2826 (.Y(N10010),.A(N9828),.B(N9827));
AND2X1 AND_tmp667 (.Y(ttmp667),.A(N8307),.B(N8269));
AND2X1 AND_tmp668 (.Y(N10013),.A(N9791),.B(ttmp667));
AND2X1 AND_tmp669 (.Y(ttmp669),.A(N8307),.B(N8269));
AND2X1 AND_tmp670 (.Y(ttmp670),.A(N9758),.B(ttmp669));
AND2X1 AND_tmp671 (.Y(N10014),.A(N9344),.B(ttmp670));
AND2X1 AND_tmp672 (.Y(ttmp672),.A(N8307),.B(N8269));
AND2X1 AND_tmp673 (.Y(ttmp673),.A(N367),.B(ttmp672));
AND2X1 AND_tmp674 (.Y(ttmp674),.A(N9754),.B(ttmp673));
AND2X1 AND_tmp675 (.Y(N10015),.A(N9344),.B(ttmp674));
AND2X1 AND_tmp676 (.Y(ttmp676),.A(N8394),.B(N8421));
AND2X1 AND_tmp677 (.Y(N10016),.A(N9786),.B(ttmp676));
AND2X1 AND_tmp678 (.Y(ttmp678),.A(N8394),.B(N8421));
AND2X1 AND_tmp679 (.Y(ttmp679),.A(N9820),.B(ttmp678));
AND2X1 AND_tmp680 (.Y(N10017),.A(N9332),.B(ttmp679));
AND2X1 AND_tmp681 (.Y(ttmp681),.A(N8394),.B(N8421));
AND2X1 AND_tmp682 (.Y(N10018),.A(N9786),.B(ttmp681));
AND2X1 AND_tmp683 (.Y(ttmp683),.A(N8394),.B(N8421));
AND2X1 AND_tmp684 (.Y(ttmp684),.A(N9820),.B(ttmp683));
AND2X1 AND_tmp685 (.Y(N10019),.A(N9332),.B(ttmp684));
AND2X1 AND_tmp686 (.Y(ttmp686),.A(N8298),.B(N8262));
AND2X1 AND_tmp687 (.Y(N10020),.A(N9809),.B(ttmp686));
AND2X1 AND_tmp688 (.Y(ttmp688),.A(N8298),.B(N8262));
AND2X1 AND_tmp689 (.Y(ttmp689),.A(N9779),.B(ttmp688));
AND2X1 AND_tmp690 (.Y(N10021),.A(N9385),.B(ttmp689));
AND2X1 AND_tmp691 (.Y(ttmp691),.A(N8298),.B(N8262));
AND2X1 AND_tmp692 (.Y(ttmp692),.A(N367),.B(ttmp691));
AND2X1 AND_tmp693 (.Y(ttmp693),.A(N9775),.B(ttmp692));
AND2X1 AND_tmp694 (.Y(N10022),.A(N9385),.B(ttmp693));
INVX1 NOT1_2837 (.Y(N10023),.A(N9945));
INVX1 NOT1_2838 (.Y(N10024),.A(N9946));
NAND2X1 NAND2_2839 (.Y(N10025),.A(N9740),.B(N9893));
INVX1 NOT1_2840 (.Y(N10026),.A(N9923));
INVX1 NOT1_2841 (.Y(N10028),.A(N9924));
NAND2X1 NAND2_2842 (.Y(N10032),.A(N8595),.B(N9897));
NAND2X1 NAND2_2843 (.Y(N10033),.A(N8598),.B(N9899));
NAND2X1 NAND2_2844 (.Y(N10034),.A(N8601),.B(N9901));
NAND2X1 NAND2_2845 (.Y(N10035),.A(N8604),.B(N9903));
NAND2X1 NAND2_2846 (.Y(N10036),.A(N4803),.B(N9906));
NAND2X1 NAND2_2847 (.Y(N10037),.A(N4806),.B(N9908));
NAND2X1 NAND2_2848 (.Y(N10038),.A(N8627),.B(N9910));
AND2X1 AND2_2849 (.Y(N10039),.A(N9809),.B(N8298));
AND2X1 AND_tmp695 (.Y(ttmp695),.A(N9385),.B(N8298));
AND2X1 AND_tmp696 (.Y(N10040),.A(N9779),.B(ttmp695));
AND2X1 AND_tmp697 (.Y(ttmp697),.A(N9385),.B(N8298));
AND2X1 AND_tmp698 (.Y(ttmp698),.A(N367),.B(ttmp697));
AND2X1 AND_tmp699 (.Y(N10041),.A(N9775),.B(ttmp698));
AND2X1 AND2_2852 (.Y(N10042),.A(N9779),.B(N9385));
AND2X1 AND_tmp700 (.Y(ttmp700),.A(N9775),.B(N9385));
AND2X1 AND_tmp701 (.Y(N10043),.A(N367),.B(ttmp700));
NAND2X1 NAND2_2854 (.Y(N10050),.A(N8727),.B(N9938));
INVX1 NOT1_2855 (.Y(N10053),.A(N9817));
AND2X1 AND2_2856 (.Y(N10054),.A(N9817),.B(N9029));
AND2X1 AND2_2857 (.Y(N10055),.A(N9786),.B(N8394));
AND2X1 AND_tmp702 (.Y(ttmp702),.A(N9332),.B(N8394));
AND2X1 AND_tmp703 (.Y(N10056),.A(N9820),.B(ttmp702));
AND2X1 AND2_2859 (.Y(N10057),.A(N9791),.B(N8307));
AND2X1 AND_tmp704 (.Y(ttmp704),.A(N9344),.B(N8307));
AND2X1 AND_tmp705 (.Y(N10058),.A(N9758),.B(ttmp704));
AND2X1 AND_tmp706 (.Y(ttmp706),.A(N9344),.B(N8307));
AND2X1 AND_tmp707 (.Y(ttmp707),.A(N367),.B(ttmp706));
AND2X1 AND_tmp708 (.Y(N10059),.A(N9754),.B(ttmp707));
AND2X1 AND2_2862 (.Y(N10060),.A(N9758),.B(N9344));
AND2X1 AND_tmp709 (.Y(ttmp709),.A(N9754),.B(N9344));
AND2X1 AND_tmp710 (.Y(N10061),.A(N367),.B(ttmp709));
NAND2X1 NAND2_2864 (.Y(N10062),.A(N4997),.B(N9947));
NAND2X1 NAND2_2865 (.Y(N10067),.A(N8811),.B(N9953));
NAND2X1 NAND2_2866 (.Y(N10070),.A(N9955),.B(N9836));
NAND2X1 NAND2_2867 (.Y(N10073),.A(N9956),.B(N9838));
NAND2X1 NAND2_2868 (.Y(N10076),.A(N9068),.B(N9957));
NAND2X1 NAND2_2869 (.Y(N10077),.A(N9074),.B(N9959));
NAND2X1 NAND2_2870 (.Y(N10082),.A(N9089),.B(N9967));
NAND2X1 NAND2_2871 (.Y(N10083),.A(N9095),.B(N9969));
NAND2X1 NAND2_2872 (.Y(N10084),.A(N4871),.B(N9971));
NAND2X1 NAND2_2873 (.Y(N10085),.A(N6214),.B(N9973));
NAND2X1 NAND2_2874 (.Y(N10086),.A(N6217),.B(N9975));
NAND2X1 NAND2_2875 (.Y(N10093),.A(N5027),.B(N9995));
NAND2X1 NAND2_2876 (.Y(N10094),.A(N6232),.B(N9997));
OR2X1 OR_tmp711 (.Y(ttmp711),.A(N10014),.B(N10015));
OR2X1 OR_tmp712 (.Y(ttmp712),.A(N9238),.B(ttmp711));
OR2X1 OR_tmp713 (.Y(ttmp713),.A(N9732),.B(ttmp712));
OR2X1 OR_tmp714 (.Y(N10101),.A(N10013),.B(ttmp713));
OR2X1 OR_tmp715 (.Y(ttmp715),.A(N10017),.B(N9734));
OR2X1 OR_tmp716 (.Y(ttmp716),.A(N9339),.B(ttmp715));
OR2X1 OR_tmp717 (.Y(ttmp717),.A(N9526),.B(ttmp716));
OR2X1 OR_tmp718 (.Y(N10102),.A(N10016),.B(ttmp717));
OR2X1 OR_tmp719 (.Y(ttmp719),.A(N10019),.B(N9735));
OR2X1 OR_tmp720 (.Y(ttmp720),.A(N9339),.B(ttmp719));
OR2X1 OR_tmp721 (.Y(ttmp721),.A(N9531),.B(ttmp720));
OR2X1 OR_tmp722 (.Y(N10103),.A(N10018),.B(ttmp721));
OR2X1 OR_tmp723 (.Y(ttmp723),.A(N10021),.B(N10022));
OR2X1 OR_tmp724 (.Y(ttmp724),.A(N9242),.B(ttmp723));
OR2X1 OR_tmp725 (.Y(ttmp725),.A(N9736),.B(ttmp724));
OR2X1 OR_tmp726 (.Y(N10104),.A(N10020),.B(ttmp725));
AND2X1 AND2_2881 (.Y(N10105),.A(N9925),.B(N9894));
AND2X1 AND2_2882 (.Y(N10106),.A(N9925),.B(N9895));
AND2X1 AND2_2883 (.Y(N10107),.A(N9925),.B(N9896));
AND2X1 AND2_2884 (.Y(N10108),.A(N9925),.B(N8253));
NAND2X1 NAND2_2885 (.Y(N10109),.A(N10032),.B(N9898));
NAND2X1 NAND2_2886 (.Y(N10110),.A(N10033),.B(N9900));
NAND2X1 NAND2_2887 (.Y(N10111),.A(N10034),.B(N9902));
NAND2X1 NAND2_2888 (.Y(N10112),.A(N10035),.B(N9904));
NAND2X1 NAND2_2889 (.Y(N10113),.A(N10036),.B(N9907));
NAND2X1 NAND2_2890 (.Y(N10114),.A(N10037),.B(N9909));
NAND2X1 NAND2_2891 (.Y(N10115),.A(N10038),.B(N9911));
OR2X1 OR_tmp727 (.Y(ttmp727),.A(N10040),.B(N10041));
OR2X1 OR_tmp728 (.Y(ttmp728),.A(N9265),.B(ttmp727));
OR2X1 OR_tmp729 (.Y(N10116),.A(N10039),.B(ttmp728));
OR2X1 OR_tmp730 (.Y(ttmp730),.A(N10042),.B(N10043));
OR2X1 OR_tmp731 (.Y(N10119),.A(N9809),.B(ttmp730));
INVX1 NOT1_2894 (.Y(N10124),.A(N9925));
AND2X1 AND2_2895 (.Y(N10130),.A(N9768),.B(N9925));
INVX1 NOT1_2896 (.Y(N10131),.A(N9932));
INVX1 NOT1_2897 (.Y(N10132),.A(N9935));
AND2X1 AND2_2898 (.Y(N10133),.A(N9932),.B(N8920));
NAND2X1 NAND2_2899 (.Y(N10134),.A(N10050),.B(N9939));
INVX1 NOT1_2900 (.Y(N10135),.A(N9983));
NAND2X1 NAND2_2901 (.Y(N10136),.A(N9983),.B(N9324));
INVX1 NOT1_2902 (.Y(N10137),.A(N9986));
NAND2X1 NAND2_2903 (.Y(N10138),.A(N9986),.B(N9784));
AND2X1 AND2_2904 (.Y(N10139),.A(N9785),.B(N10053));
OR2X1 OR_tmp732 (.Y(ttmp732),.A(N10056),.B(N9790));
OR2X1 OR_tmp733 (.Y(ttmp733),.A(N8943),.B(ttmp732));
OR2X1 OR_tmp734 (.Y(N10140),.A(N10055),.B(ttmp733));
OR2X1 OR_tmp735 (.Y(ttmp735),.A(N10058),.B(N10059));
OR2X1 OR_tmp736 (.Y(ttmp736),.A(N9268),.B(ttmp735));
OR2X1 OR_tmp737 (.Y(N10141),.A(N10057),.B(ttmp736));
OR2X1 OR_tmp738 (.Y(ttmp738),.A(N10060),.B(N10061));
OR2X1 OR_tmp739 (.Y(N10148),.A(N9791),.B(ttmp738));
NAND2X1 NAND2_2908 (.Y(N10155),.A(N10062),.B(N9948));
INVX1 NOT1_2909 (.Y(N10156),.A(N9989));
NAND2X1 NAND2_2910 (.Y(N10157),.A(N9989),.B(N9805));
INVX1 NOT1_2911 (.Y(N10158),.A(N9992));
NAND2X1 NAND2_2912 (.Y(N10159),.A(N9992),.B(N9806));
INVX1 NOT1_2913 (.Y(N10160),.A(N9949));
NAND2X1 NAND2_2914 (.Y(N10161),.A(N10067),.B(N9954));
INVX1 NOT1_2915 (.Y(N10162),.A(N10007));
NAND2X1 NAND2_2916 (.Y(N10163),.A(N10007),.B(N9825));
INVX1 NOT1_2917 (.Y(N10164),.A(N10010));
NAND2X1 NAND2_2918 (.Y(N10165),.A(N10010),.B(N9826));
NAND2X1 NAND2_2919 (.Y(N10170),.A(N10076),.B(N9958));
NAND2X1 NAND2_2920 (.Y(N10173),.A(N10077),.B(N9960));
INVX1 NOT1_2921 (.Y(N10176),.A(N9961));
NAND2X1 NAND2_2922 (.Y(N10177),.A(N9961),.B(N9082));
INVX1 NOT1_2923 (.Y(N10178),.A(N9964));
NAND2X1 NAND2_2924 (.Y(N10179),.A(N9964),.B(N9086));
NAND2X1 NAND2_2925 (.Y(N10180),.A(N10082),.B(N9968));
NAND2X1 NAND2_2926 (.Y(N10183),.A(N10083),.B(N9970));
NAND2X1 NAND2_2927 (.Y(N10186),.A(N9972),.B(N10084));
NAND2X1 NAND2_2928 (.Y(N10189),.A(N9974),.B(N10085));
NAND2X1 NAND2_2929 (.Y(N10192),.A(N9976),.B(N10086));
INVX1 NOT1_2930 (.Y(N10195),.A(N9979));
NAND2X1 NAND2_2931 (.Y(N10196),.A(N9979),.B(N9982));
NAND2X1 NAND2_2932 (.Y(N10197),.A(N9996),.B(N10093));
NAND2X1 NAND2_2933 (.Y(N10200),.A(N9998),.B(N10094));
INVX1 NOT1_2934 (.Y(N10203),.A(N9999));
NAND2X1 NAND2_2935 (.Y(N10204),.A(N9999),.B(N10002));
INVX1 NOT1_2936 (.Y(N10205),.A(N10003));
NAND2X1 NAND2_2937 (.Y(N10206),.A(N10003),.B(N10006));
NAND2X1 NAND2_2938 (.Y(N10212),.A(N10070),.B(N4308));
NAND2X1 NAND2_2939 (.Y(N10213),.A(N10073),.B(N4313));
AND2X1 AND2_2940 (.Y(N10230),.A(N9774),.B(N10131));
NAND2X1 NAND2_2941 (.Y(N10231),.A(N8730),.B(N10135));
NAND2X1 NAND2_2942 (.Y(N10232),.A(N9478),.B(N10137));
OR2X1 OR2_2943 (.Y(N10233),.A(N10139),.B(N10054));
NAND2X1 NAND2_2944 (.Y(N10234),.A(N7100),.B(N10140));
NAND2X1 NAND2_2945 (.Y(N10237),.A(N9485),.B(N10156));
NAND2X1 NAND2_2946 (.Y(N10238),.A(N9488),.B(N10158));
NAND2X1 NAND2_2947 (.Y(N10239),.A(N9517),.B(N10162));
NAND2X1 NAND2_2948 (.Y(N10240),.A(N9520),.B(N10164));
INVX1 NOT1_2949 (.Y(N10241),.A(N10070));
INVX1 NOT1_2950 (.Y(N10242),.A(N10073));
NAND2X1 NAND2_2951 (.Y(N10247),.A(N8146),.B(N10176));
NAND2X1 NAND2_2952 (.Y(N10248),.A(N8156),.B(N10178));
NAND2X1 NAND2_2953 (.Y(N10259),.A(N9692),.B(N10195));
NAND2X1 NAND2_2954 (.Y(N10264),.A(N9717),.B(N10203));
NAND2X1 NAND2_2955 (.Y(N10265),.A(N9723),.B(N10205));
AND2X1 AND2_2956 (.Y(N10266),.A(N10026),.B(N10124));
AND2X1 AND2_2957 (.Y(N10267),.A(N10028),.B(N10124));
AND2X1 AND2_2958 (.Y(N10268),.A(N9742),.B(N10124));
AND2X1 AND2_2959 (.Y(N10269),.A(N6923),.B(N10124));
NAND2X1 NAND2_2960 (.Y(N10270),.A(N6762),.B(N10116));
NAND2X1 NAND2_2961 (.Y(N10271),.A(N3061),.B(N10241));
NAND2X1 NAND2_2962 (.Y(N10272),.A(N3064),.B(N10242));
BUFX1 BUFF1_2963 (.Y(N10273),.A(N10116));
AND2X1 AND_tmp740 (.Y(ttmp740),.A(N5718),.B(N5697));
AND2X1 AND_tmp741 (.Y(ttmp741),.A(N10141),.B(ttmp740));
AND2X1 AND_tmp742 (.Y(ttmp742),.A(N5728),.B(ttmp741));
AND2X1 AND_tmp743 (.Y(N10278),.A(N5707),.B(ttmp742));
AND2X1 AND_tmp744 (.Y(ttmp744),.A(N5707),.B(N5718));
AND2X1 AND_tmp745 (.Y(ttmp745),.A(N10141),.B(ttmp744));
AND2X1 AND_tmp746 (.Y(N10279),.A(N5728),.B(ttmp745));
AND2X1 AND_tmp747 (.Y(ttmp747),.A(N5728),.B(N5718));
AND2X1 AND_tmp748 (.Y(N10280),.A(N10141),.B(ttmp747));
AND2X1 AND2_2967 (.Y(N10281),.A(N10141),.B(N5728));
AND2X1 AND2_2968 (.Y(N10282),.A(N6784),.B(N10141));
INVX1 NOT1_2969 (.Y(N10283),.A(N10119));
AND2X1 AND_tmp749 (.Y(ttmp749),.A(N5926),.B(N5905));
AND2X1 AND_tmp750 (.Y(ttmp750),.A(N10148),.B(ttmp749));
AND2X1 AND_tmp751 (.Y(ttmp751),.A(N5936),.B(ttmp750));
AND2X1 AND_tmp752 (.Y(N10287),.A(N5915),.B(ttmp751));
AND2X1 AND_tmp753 (.Y(ttmp753),.A(N5915),.B(N5926));
AND2X1 AND_tmp754 (.Y(ttmp754),.A(N10148),.B(ttmp753));
AND2X1 AND_tmp755 (.Y(N10288),.A(N5936),.B(ttmp754));
AND2X1 AND_tmp756 (.Y(ttmp756),.A(N5936),.B(N5926));
AND2X1 AND_tmp757 (.Y(N10289),.A(N10148),.B(ttmp756));
AND2X1 AND2_2973 (.Y(N10290),.A(N10148),.B(N5936));
AND2X1 AND2_2974 (.Y(N10291),.A(N6881),.B(N10148));
AND2X1 AND2_2975 (.Y(N10292),.A(N8898),.B(N10124));
NAND2X1 NAND2_2976 (.Y(N10293),.A(N10231),.B(N10136));
NAND2X1 NAND2_2977 (.Y(N10294),.A(N10232),.B(N10138));
NAND2X1 NAND2_2978 (.Y(N10295),.A(N8412),.B(N10233));
AND2X1 AND2_2979 (.Y(N10296),.A(N8959),.B(N10234));
NAND2X1 NAND2_2980 (.Y(N10299),.A(N10237),.B(N10157));
NAND2X1 NAND2_2981 (.Y(N10300),.A(N10238),.B(N10159));
OR2X1 OR2_2982 (.Y(N10301),.A(N10230),.B(N10133));
NAND2X1 NAND2_2983 (.Y(N10306),.A(N10239),.B(N10163));
NAND2X1 NAND2_2984 (.Y(N10307),.A(N10240),.B(N10165));
BUFX1 BUFF1_2985 (.Y(N10308),.A(N10148));
BUFX1 BUFF1_2986 (.Y(N10311),.A(N10141));
INVX1 NOT1_2987 (.Y(N10314),.A(N10170));
NAND2X1 NAND2_2988 (.Y(N10315),.A(N10170),.B(N9071));
INVX1 NOT1_2989 (.Y(N10316),.A(N10173));
NAND2X1 NAND2_2990 (.Y(N10317),.A(N10173),.B(N9077));
NAND2X1 NAND2_2991 (.Y(N10318),.A(N10247),.B(N10177));
NAND2X1 NAND2_2992 (.Y(N10321),.A(N10248),.B(N10179));
INVX1 NOT1_2993 (.Y(N10324),.A(N10180));
NAND2X1 NAND2_2994 (.Y(N10325),.A(N10180),.B(N9092));
INVX1 NOT1_2995 (.Y(N10326),.A(N10183));
NAND2X1 NAND2_2996 (.Y(N10327),.A(N10183),.B(N9098));
INVX1 NOT1_2997 (.Y(N10328),.A(N10186));
NAND2X1 NAND2_2998 (.Y(N10329),.A(N10186),.B(N9674));
INVX1 NOT1_2999 (.Y(N10330),.A(N10189));
NAND2X1 NAND2_3000 (.Y(N10331),.A(N10189),.B(N9678));
INVX1 NOT1_3001 (.Y(N10332),.A(N10192));
NAND2X1 NAND2_3002 (.Y(N10333),.A(N10192),.B(N9977));
NAND2X1 NAND2_3003 (.Y(N10334),.A(N10259),.B(N10196));
INVX1 NOT1_3004 (.Y(N10337),.A(N10197));
NAND2X1 NAND2_3005 (.Y(N10338),.A(N10197),.B(N9710));
INVX1 NOT1_3006 (.Y(N10339),.A(N10200));
NAND2X1 NAND2_3007 (.Y(N10340),.A(N10200),.B(N9714));
NAND2X1 NAND2_3008 (.Y(N10341),.A(N10264),.B(N10204));
NAND2X1 NAND2_3009 (.Y(N10344),.A(N10265),.B(N10206));
OR2X1 OR2_3010 (.Y(N10350),.A(N10266),.B(N10105));
OR2X1 OR2_3011 (.Y(N10351),.A(N10267),.B(N10106));
OR2X1 OR2_3012 (.Y(N10352),.A(N10268),.B(N10107));
OR2X1 OR2_3013 (.Y(N10353),.A(N10269),.B(N10108));
AND2X1 AND2_3014 (.Y(N10354),.A(N8857),.B(N10270));
NAND2X1 NAND2_3015 (.Y(N10357),.A(N10271),.B(N10212));
NAND2X1 NAND2_3016 (.Y(N10360),.A(N10272),.B(N10213));
OR2X1 OR2_3017 (.Y(N10367),.A(N7620),.B(N10282));
OR2X1 OR2_3018 (.Y(N10375),.A(N7671),.B(N10291));
OR2X1 OR2_3019 (.Y(N10381),.A(N10292),.B(N10130));
AND2X1 AND_tmp758 (.Y(ttmp758),.A(N10293),.B(N10294));
AND2X1 AND_tmp759 (.Y(ttmp759),.A(N10114),.B(ttmp758));
AND2X1 AND_tmp760 (.Y(N10388),.A(N10134),.B(ttmp759));
AND2X1 AND2_3021 (.Y(N10391),.A(N9582),.B(N10295));
AND2X1 AND_tmp761 (.Y(ttmp761),.A(N10299),.B(N10300));
AND2X1 AND_tmp762 (.Y(ttmp762),.A(N10113),.B(ttmp761));
AND2X1 AND_tmp763 (.Y(N10399),.A(N10115),.B(ttmp762));
AND2X1 AND_tmp764 (.Y(ttmp764),.A(N10306),.B(N10307));
AND2X1 AND_tmp765 (.Y(ttmp765),.A(N10155),.B(ttmp764));
AND2X1 AND_tmp766 (.Y(N10402),.A(N10161),.B(ttmp765));
OR2X1 OR_tmp767 (.Y(ttmp767),.A(N6890),.B(N10287));
OR2X1 OR_tmp768 (.Y(ttmp768),.A(N3229),.B(ttmp767));
OR2X1 OR_tmp769 (.Y(ttmp769),.A(N6888),.B(ttmp768));
OR2X1 OR_tmp770 (.Y(N10406),.A(N6889),.B(ttmp769));
OR2X1 OR_tmp771 (.Y(ttmp771),.A(N6892),.B(N10288));
OR2X1 OR_tmp772 (.Y(ttmp772),.A(N3232),.B(ttmp771));
OR2X1 OR_tmp773 (.Y(N10409),.A(N6891),.B(ttmp772));
OR2X1 OR_tmp774 (.Y(ttmp774),.A(N6893),.B(N10289));
OR2X1 OR_tmp775 (.Y(N10412),.A(N3236),.B(ttmp774));
OR2X1 OR2_3027 (.Y(N10415),.A(N3241),.B(N10290));
OR2X1 OR_tmp776 (.Y(ttmp776),.A(N6793),.B(N10278));
OR2X1 OR_tmp777 (.Y(ttmp777),.A(N3137),.B(ttmp776));
OR2X1 OR_tmp778 (.Y(ttmp778),.A(N6791),.B(ttmp777));
OR2X1 OR_tmp779 (.Y(N10419),.A(N6792),.B(ttmp778));
OR2X1 OR_tmp780 (.Y(ttmp780),.A(N6795),.B(N10279));
OR2X1 OR_tmp781 (.Y(ttmp781),.A(N3140),.B(ttmp780));
OR2X1 OR_tmp782 (.Y(N10422),.A(N6794),.B(ttmp781));
OR2X1 OR_tmp783 (.Y(ttmp783),.A(N6796),.B(N10280));
OR2X1 OR_tmp784 (.Y(N10425),.A(N3144),.B(ttmp783));
OR2X1 OR2_3031 (.Y(N10428),.A(N3149),.B(N10281));
NAND2X1 NAND2_3032 (.Y(N10431),.A(N8117),.B(N10314));
NAND2X1 NAND2_3033 (.Y(N10432),.A(N8134),.B(N10316));
NAND2X1 NAND2_3034 (.Y(N10437),.A(N8169),.B(N10324));
NAND2X1 NAND2_3035 (.Y(N10438),.A(N8186),.B(N10326));
NAND2X1 NAND2_3036 (.Y(N10439),.A(N9117),.B(N10328));
NAND2X1 NAND2_3037 (.Y(N10440),.A(N9127),.B(N10330));
NAND2X1 NAND2_3038 (.Y(N10441),.A(N9682),.B(N10332));
NAND2X1 NAND2_3039 (.Y(N10444),.A(N9183),.B(N10337));
NAND2X1 NAND2_3040 (.Y(N10445),.A(N9193),.B(N10339));
INVX1 NOT1_3041 (.Y(N10450),.A(N10296));
AND2X1 AND2_3042 (.Y(N10451),.A(N10296),.B(N4193));
INVX1 NOT1_3043 (.Y(N10455),.A(N10308));
NAND2X1 NAND2_3044 (.Y(N10456),.A(N10308),.B(N8242));
INVX1 NOT1_3045 (.Y(N10465),.A(N10311));
NAND2X1 NAND2_3046 (.Y(N10466),.A(N10311),.B(N8247));
INVX1 NOT1_3047 (.Y(N10479),.A(N10273));
INVX1 NOT1_3048 (.Y(N10497),.A(N10301));
NAND2X1 NAND2_3049 (.Y(N10509),.A(N10431),.B(N10315));
NAND2X1 NAND2_3050 (.Y(N10512),.A(N10432),.B(N10317));
INVX1 NOT1_3051 (.Y(N10515),.A(N10318));
NAND2X1 NAND2_3052 (.Y(N10516),.A(N10318),.B(N8632));
INVX1 NOT1_3053 (.Y(N10517),.A(N10321));
NAND2X1 NAND2_3054 (.Y(N10518),.A(N10321),.B(N8637));
NAND2X1 NAND2_3055 (.Y(N10519),.A(N10437),.B(N10325));
NAND2X1 NAND2_3056 (.Y(N10522),.A(N10438),.B(N10327));
NAND2X1 NAND2_3057 (.Y(N10525),.A(N10439),.B(N10329));
NAND2X1 NAND2_3058 (.Y(N10528),.A(N10440),.B(N10331));
NAND2X1 NAND2_3059 (.Y(N10531),.A(N10441),.B(N10333));
INVX1 NOT1_3060 (.Y(N10534),.A(N10334));
NAND2X1 NAND2_3061 (.Y(N10535),.A(N10334),.B(N9695));
NAND2X1 NAND2_3062 (.Y(N10536),.A(N10444),.B(N10338));
NAND2X1 NAND2_3063 (.Y(N10539),.A(N10445),.B(N10340));
INVX1 NOT1_3064 (.Y(N10542),.A(N10341));
NAND2X1 NAND2_3065 (.Y(N10543),.A(N10341),.B(N9720));
INVX1 NOT1_3066 (.Y(N10544),.A(N10344));
NAND2X1 NAND2_3067 (.Y(N10545),.A(N10344),.B(N9726));
AND2X1 AND2_3068 (.Y(N10546),.A(N5631),.B(N10450));
INVX1 NOT1_3069 (.Y(N10547),.A(N10391));
AND2X1 AND2_3070 (.Y(N10548),.A(N10391),.B(N8950));
AND2X1 AND2_3071 (.Y(N10549),.A(N5165),.B(N10367));
INVX1 NOT1_3072 (.Y(N10550),.A(N10354));
AND2X1 AND2_3073 (.Y(N10551),.A(N10354),.B(N3126));
NAND2X1 NAND2_3074 (.Y(N10552),.A(N7411),.B(N10455));
AND2X1 AND2_3075 (.Y(N10553),.A(N10375),.B(N9539));
AND2X1 AND2_3076 (.Y(N10554),.A(N10375),.B(N9540));
AND2X1 AND2_3077 (.Y(N10555),.A(N10375),.B(N9541));
AND2X1 AND2_3078 (.Y(N10556),.A(N10375),.B(N6761));
INVX1 NOT1_3079 (.Y(N10557),.A(N10406));
NAND2X1 NAND2_3080 (.Y(N10558),.A(N10406),.B(N8243));
INVX1 NOT1_3081 (.Y(N10559),.A(N10409));
NAND2X1 NAND2_3082 (.Y(N10560),.A(N10409),.B(N8244));
INVX1 NOT1_3083 (.Y(N10561),.A(N10412));
NAND2X1 NAND2_3084 (.Y(N10562),.A(N10412),.B(N8245));
INVX1 NOT1_3085 (.Y(N10563),.A(N10415));
NAND2X1 NAND2_3086 (.Y(N10564),.A(N10415),.B(N8246));
NAND2X1 NAND2_3087 (.Y(N10565),.A(N7426),.B(N10465));
INVX1 NOT1_3088 (.Y(N10566),.A(N10419));
NAND2X1 NAND2_3089 (.Y(N10567),.A(N10419),.B(N8248));
INVX1 NOT1_3090 (.Y(N10568),.A(N10422));
NAND2X1 NAND2_3091 (.Y(N10569),.A(N10422),.B(N8249));
INVX1 NOT1_3092 (.Y(N10570),.A(N10425));
NAND2X1 NAND2_3093 (.Y(N10571),.A(N10425),.B(N8250));
INVX1 NOT1_3094 (.Y(N10572),.A(N10428));
NAND2X1 NAND2_3095 (.Y(N10573),.A(N10428),.B(N8251));
INVX1 NOT1_3096 (.Y(N10574),.A(N10399));
INVX1 NOT1_3097 (.Y(N10575),.A(N10402));
INVX1 NOT1_3098 (.Y(N10576),.A(N10388));
AND2X1 AND_tmp785 (.Y(ttmp785),.A(N10402),.B(N10388));
AND2X1 AND_tmp786 (.Y(N10577),.A(N10399),.B(ttmp785));
AND2X1 AND_tmp787 (.Y(ttmp787),.A(N9543),.B(N10273));
AND2X1 AND_tmp788 (.Y(N10581),.A(N10360),.B(ttmp787));
AND2X1 AND_tmp789 (.Y(ttmp789),.A(N9905),.B(N10273));
AND2X1 AND_tmp790 (.Y(N10582),.A(N10357),.B(ttmp789));
INVX1 NOT1_3102 (.Y(N10583),.A(N10367));
AND2X1 AND2_3103 (.Y(N10587),.A(N10367),.B(N5735));
AND2X1 AND2_3104 (.Y(N10588),.A(N10367),.B(N3135));
INVX1 NOT1_3105 (.Y(N10589),.A(N10375));
AND2X1 AND_tmp791 (.Y(ttmp791),.A(N7170),.B(N7149));
AND2X1 AND_tmp792 (.Y(ttmp792),.A(N10381),.B(ttmp791));
AND2X1 AND_tmp793 (.Y(ttmp793),.A(N7180),.B(ttmp792));
AND2X1 AND_tmp794 (.Y(N10594),.A(N7159),.B(ttmp793));
AND2X1 AND_tmp795 (.Y(ttmp795),.A(N7159),.B(N7170));
AND2X1 AND_tmp796 (.Y(ttmp796),.A(N10381),.B(ttmp795));
AND2X1 AND_tmp797 (.Y(N10595),.A(N7180),.B(ttmp796));
AND2X1 AND_tmp798 (.Y(ttmp798),.A(N7180),.B(N7170));
AND2X1 AND_tmp799 (.Y(N10596),.A(N10381),.B(ttmp798));
AND2X1 AND2_3109 (.Y(N10597),.A(N10381),.B(N7180));
AND2X1 AND2_3110 (.Y(N10598),.A(N8444),.B(N10381));
BUFX1 BUFF1_3111 (.Y(N10602),.A(N10381));
NAND2X1 NAND2_3112 (.Y(N10609),.A(N7479),.B(N10515));
NAND2X1 NAND2_3113 (.Y(N10610),.A(N7491),.B(N10517));
NAND2X1 NAND2_3114 (.Y(N10621),.A(N9149),.B(N10534));
NAND2X1 NAND2_3115 (.Y(N10626),.A(N9206),.B(N10542));
NAND2X1 NAND2_3116 (.Y(N10627),.A(N9223),.B(N10544));
OR2X1 OR2_3117 (.Y(N10628),.A(N10546),.B(N10451));
AND2X1 AND2_3118 (.Y(N10629),.A(N9733),.B(N10547));
AND2X1 AND2_3119 (.Y(N10631),.A(N5166),.B(N10550));
NAND2X1 NAND2_3120 (.Y(N10632),.A(N10552),.B(N10456));
NAND2X1 NAND2_3121 (.Y(N10637),.A(N7414),.B(N10557));
NAND2X1 NAND2_3122 (.Y(N10638),.A(N7417),.B(N10559));
NAND2X1 NAND2_3123 (.Y(N10639),.A(N7420),.B(N10561));
NAND2X1 NAND2_3124 (.Y(N10640),.A(N7423),.B(N10563));
NAND2X1 NAND2_3125 (.Y(N10641),.A(N10565),.B(N10466));
NAND2X1 NAND2_3126 (.Y(N10642),.A(N7429),.B(N10566));
NAND2X1 NAND2_3127 (.Y(N10643),.A(N7432),.B(N10568));
NAND2X1 NAND2_3128 (.Y(N10644),.A(N7435),.B(N10570));
NAND2X1 NAND2_3129 (.Y(N10645),.A(N7438),.B(N10572));
AND2X1 AND_tmp800 (.Y(ttmp800),.A(N887),.B(N10577));
AND2X1 AND_tmp801 (.Y(N10647),.A(N886),.B(ttmp800));
AND2X1 AND_tmp802 (.Y(ttmp802),.A(N8857),.B(N10479));
AND2X1 AND_tmp803 (.Y(N10648),.A(N10360),.B(ttmp802));
AND2X1 AND_tmp804 (.Y(ttmp804),.A(N7609),.B(N10479));
AND2X1 AND_tmp805 (.Y(N10649),.A(N10357),.B(ttmp804));
OR2X1 OR2_3133 (.Y(N10652),.A(N8966),.B(N10598));
OR2X1 OR_tmp806 (.Y(ttmp806),.A(N8453),.B(N10594));
OR2X1 OR_tmp807 (.Y(ttmp807),.A(N4675),.B(ttmp806));
OR2X1 OR_tmp808 (.Y(ttmp808),.A(N8451),.B(ttmp807));
OR2X1 OR_tmp809 (.Y(N10659),.A(N8452),.B(ttmp808));
OR2X1 OR_tmp810 (.Y(ttmp810),.A(N8455),.B(N10595));
OR2X1 OR_tmp811 (.Y(ttmp811),.A(N4678),.B(ttmp810));
OR2X1 OR_tmp812 (.Y(N10662),.A(N8454),.B(ttmp811));
OR2X1 OR_tmp813 (.Y(ttmp813),.A(N8456),.B(N10596));
OR2X1 OR_tmp814 (.Y(N10665),.A(N4682),.B(ttmp813));
OR2X1 OR2_3137 (.Y(N10668),.A(N4687),.B(N10597));
INVX1 NOT1_3138 (.Y(N10671),.A(N10509));
NAND2X1 NAND2_3139 (.Y(N10672),.A(N10509),.B(N8615));
INVX1 NOT1_3140 (.Y(N10673),.A(N10512));
NAND2X1 NAND2_3141 (.Y(N10674),.A(N10512),.B(N8624));
NAND2X1 NAND2_3142 (.Y(N10675),.A(N10609),.B(N10516));
NAND2X1 NAND2_3143 (.Y(N10678),.A(N10610),.B(N10518));
INVX1 NOT1_3144 (.Y(N10681),.A(N10519));
NAND2X1 NAND2_3145 (.Y(N10682),.A(N10519),.B(N8644));
INVX1 NOT1_3146 (.Y(N10683),.A(N10522));
NAND2X1 NAND2_3147 (.Y(N10684),.A(N10522),.B(N8653));
INVX1 NOT1_3148 (.Y(N10685),.A(N10525));
NAND2X1 NAND2_3149 (.Y(N10686),.A(N10525),.B(N9454));
INVX1 NOT1_3150 (.Y(N10687),.A(N10528));
NAND2X1 NAND2_3151 (.Y(N10688),.A(N10528),.B(N9459));
INVX1 NOT1_3152 (.Y(N10689),.A(N10531));
NAND2X1 NAND2_3153 (.Y(N10690),.A(N10531),.B(N9978));
NAND2X1 NAND2_3154 (.Y(N10691),.A(N10621),.B(N10535));
INVX1 NOT1_3155 (.Y(N10694),.A(N10536));
NAND2X1 NAND2_3156 (.Y(N10695),.A(N10536),.B(N9493));
INVX1 NOT1_3157 (.Y(N10696),.A(N10539));
NAND2X1 NAND2_3158 (.Y(N10697),.A(N10539),.B(N9498));
NAND2X1 NAND2_3159 (.Y(N10698),.A(N10626),.B(N10543));
NAND2X1 NAND2_3160 (.Y(N10701),.A(N10627),.B(N10545));
OR2X1 OR2_3161 (.Y(N10704),.A(N10629),.B(N10548));
AND2X1 AND2_3162 (.Y(N10705),.A(N3159),.B(N10583));
OR2X1 OR2_3163 (.Y(N10706),.A(N10631),.B(N10551));
AND2X1 AND2_3164 (.Y(N10707),.A(N9737),.B(N10589));
AND2X1 AND2_3165 (.Y(N10708),.A(N9738),.B(N10589));
AND2X1 AND2_3166 (.Y(N10709),.A(N9243),.B(N10589));
AND2X1 AND2_3167 (.Y(N10710),.A(N5892),.B(N10589));
NAND2X1 NAND2_3168 (.Y(N10711),.A(N10637),.B(N10558));
NAND2X1 NAND2_3169 (.Y(N10712),.A(N10638),.B(N10560));
NAND2X1 NAND2_3170 (.Y(N10713),.A(N10639),.B(N10562));
NAND2X1 NAND2_3171 (.Y(N10714),.A(N10640),.B(N10564));
NAND2X1 NAND2_3172 (.Y(N10715),.A(N10642),.B(N10567));
NAND2X1 NAND2_3173 (.Y(N10716),.A(N10643),.B(N10569));
NAND2X1 NAND2_3174 (.Y(N10717),.A(N10644),.B(N10571));
NAND2X1 NAND2_3175 (.Y(N10718),.A(N10645),.B(N10573));
INVX1 NOT1_3176 (.Y(N10719),.A(N10602));
NAND2X1 NAND2_3177 (.Y(N10720),.A(N10602),.B(N9244));
INVX1 NOT1_3178 (.Y(N10729),.A(N10647));
AND2X1 AND2_3179 (.Y(N10730),.A(N5178),.B(N10583));
AND2X1 AND2_3180 (.Y(N10731),.A(N2533),.B(N10583));
NAND2X1 NAND2_3181 (.Y(N10737),.A(N7447),.B(N10671));
NAND2X1 NAND2_3182 (.Y(N10738),.A(N7465),.B(N10673));
OR2X1 OR_tmp815 (.Y(ttmp815),.A(N10581),.B(N10582));
OR2X1 OR_tmp816 (.Y(ttmp816),.A(N10648),.B(ttmp815));
OR2X1 OR_tmp817 (.Y(N10739),.A(N10649),.B(ttmp816));
NAND2X1 NAND2_3184 (.Y(N10746),.A(N7503),.B(N10681));
NAND2X1 NAND2_3185 (.Y(N10747),.A(N7521),.B(N10683));
NAND2X1 NAND2_3186 (.Y(N10748),.A(N8678),.B(N10685));
NAND2X1 NAND2_3187 (.Y(N10749),.A(N8690),.B(N10687));
NAND2X1 NAND2_3188 (.Y(N10750),.A(N9685),.B(N10689));
NAND2X1 NAND2_3189 (.Y(N10753),.A(N8757),.B(N10694));
NAND2X1 NAND2_3190 (.Y(N10754),.A(N8769),.B(N10696));
OR2X1 OR2_3191 (.Y(N10759),.A(N10705),.B(N10549));
OR2X1 OR2_3192 (.Y(N10760),.A(N10707),.B(N10553));
OR2X1 OR2_3193 (.Y(N10761),.A(N10708),.B(N10554));
OR2X1 OR2_3194 (.Y(N10762),.A(N10709),.B(N10555));
OR2X1 OR2_3195 (.Y(N10763),.A(N10710),.B(N10556));
NAND2X1 NAND2_3196 (.Y(N10764),.A(N8580),.B(N10719));
AND2X1 AND2_3197 (.Y(N10765),.A(N10652),.B(N9890));
AND2X1 AND2_3198 (.Y(N10766),.A(N10652),.B(N9891));
AND2X1 AND2_3199 (.Y(N10767),.A(N10652),.B(N9892));
AND2X1 AND2_3200 (.Y(N10768),.A(N10652),.B(N8252));
INVX1 NOT1_3201 (.Y(N10769),.A(N10659));
NAND2X1 NAND2_3202 (.Y(N10770),.A(N10659),.B(N9245));
INVX1 NOT1_3203 (.Y(N10771),.A(N10662));
NAND2X1 NAND2_3204 (.Y(N10772),.A(N10662),.B(N9246));
INVX1 NOT1_3205 (.Y(N10773),.A(N10665));
NAND2X1 NAND2_3206 (.Y(N10774),.A(N10665),.B(N9247));
INVX1 NOT1_3207 (.Y(N10775),.A(N10668));
NAND2X1 NAND2_3208 (.Y(N10776),.A(N10668),.B(N9248));
OR2X1 OR2_3209 (.Y(N10778),.A(N10730),.B(N10587));
OR2X1 OR2_3210 (.Y(N10781),.A(N10731),.B(N10588));
INVX1 NOT1_3211 (.Y(N10784),.A(N10652));
NAND2X1 NAND2_3212 (.Y(N10789),.A(N10737),.B(N10672));
NAND2X1 NAND2_3213 (.Y(N10792),.A(N10738),.B(N10674));
INVX1 NOT1_3214 (.Y(N10796),.A(N10675));
NAND2X1 NAND2_3215 (.Y(N10797),.A(N10675),.B(N8633));
INVX1 NOT1_3216 (.Y(N10798),.A(N10678));
NAND2X1 NAND2_3217 (.Y(N10799),.A(N10678),.B(N8638));
NAND2X1 NAND2_3218 (.Y(N10800),.A(N10746),.B(N10682));
NAND2X1 NAND2_3219 (.Y(N10803),.A(N10747),.B(N10684));
NAND2X1 NAND2_3220 (.Y(N10806),.A(N10748),.B(N10686));
NAND2X1 NAND2_3221 (.Y(N10809),.A(N10749),.B(N10688));
NAND2X1 NAND2_3222 (.Y(N10812),.A(N10750),.B(N10690));
INVX1 NOT1_3223 (.Y(N10815),.A(N10691));
NAND2X1 NAND2_3224 (.Y(N10816),.A(N10691),.B(N9866));
NAND2X1 NAND2_3225 (.Y(N10817),.A(N10753),.B(N10695));
NAND2X1 NAND2_3226 (.Y(N10820),.A(N10754),.B(N10697));
INVX1 NOT1_3227 (.Y(N10823),.A(N10698));
NAND2X1 NAND2_3228 (.Y(N10824),.A(N10698),.B(N9505));
INVX1 NOT1_3229 (.Y(N10825),.A(N10701));
NAND2X1 NAND2_3230 (.Y(N10826),.A(N10701),.B(N9514));
NAND2X1 NAND2_3231 (.Y(N10827),.A(N10764),.B(N10720));
NAND2X1 NAND2_3232 (.Y(N10832),.A(N8583),.B(N10769));
NAND2X1 NAND2_3233 (.Y(N10833),.A(N8586),.B(N10771));
NAND2X1 NAND2_3234 (.Y(N10834),.A(N8589),.B(N10773));
NAND2X1 NAND2_3235 (.Y(N10835),.A(N8592),.B(N10775));
INVX1 NOT1_3236 (.Y(N10836),.A(N10739));
BUFX1 BUFF1_3237 (.Y(N10837),.A(N10778));
BUFX1 BUFF1_3238 (.Y(N10838),.A(N10778));
BUFX1 BUFF1_3239 (.Y(N10839),.A(N10781));
BUFX1 BUFF1_3240 (.Y(N10840),.A(N10781));
NAND2X1 NAND2_3241 (.Y(N10845),.A(N7482),.B(N10796));
NAND2X1 NAND2_3242 (.Y(N10846),.A(N7494),.B(N10798));
NAND2X1 NAND2_3243 (.Y(N10857),.A(N9473),.B(N10815));
NAND2X1 NAND2_3244 (.Y(N10862),.A(N8781),.B(N10823));
NAND2X1 NAND2_3245 (.Y(N10863),.A(N8799),.B(N10825));
AND2X1 AND2_3246 (.Y(N10864),.A(N10023),.B(N10784));
AND2X1 AND2_3247 (.Y(N10865),.A(N10024),.B(N10784));
AND2X1 AND2_3248 (.Y(N10866),.A(N9739),.B(N10784));
AND2X1 AND2_3249 (.Y(N10867),.A(N7136),.B(N10784));
NAND2X1 NAND2_3250 (.Y(N10868),.A(N10832),.B(N10770));
NAND2X1 NAND2_3251 (.Y(N10869),.A(N10833),.B(N10772));
NAND2X1 NAND2_3252 (.Y(N10870),.A(N10834),.B(N10774));
NAND2X1 NAND2_3253 (.Y(N10871),.A(N10835),.B(N10776));
INVX1 NOT1_3254 (.Y(N10872),.A(N10789));
NAND2X1 NAND2_3255 (.Y(N10873),.A(N10789),.B(N8616));
INVX1 NOT1_3256 (.Y(N10874),.A(N10792));
NAND2X1 NAND2_3257 (.Y(N10875),.A(N10792),.B(N8625));
NAND2X1 NAND2_3258 (.Y(N10876),.A(N10845),.B(N10797));
NAND2X1 NAND2_3259 (.Y(N10879),.A(N10846),.B(N10799));
INVX1 NOT1_3260 (.Y(N10882),.A(N10800));
NAND2X1 NAND2_3261 (.Y(N10883),.A(N10800),.B(N8645));
INVX1 NOT1_3262 (.Y(N10884),.A(N10803));
NAND2X1 NAND2_3263 (.Y(N10885),.A(N10803),.B(N8654));
INVX1 NOT1_3264 (.Y(N10886),.A(N10806));
NAND2X1 NAND2_3265 (.Y(N10887),.A(N10806),.B(N9455));
INVX1 NOT1_3266 (.Y(N10888),.A(N10809));
NAND2X1 NAND2_3267 (.Y(N10889),.A(N10809),.B(N9460));
INVX1 NOT1_3268 (.Y(N10890),.A(N10812));
NAND2X1 NAND2_3269 (.Y(N10891),.A(N10812),.B(N9862));
NAND2X1 NAND2_3270 (.Y(N10892),.A(N10857),.B(N10816));
INVX1 NOT1_3271 (.Y(N10895),.A(N10817));
NAND2X1 NAND2_3272 (.Y(N10896),.A(N10817),.B(N9494));
INVX1 NOT1_3273 (.Y(N10897),.A(N10820));
NAND2X1 NAND2_3274 (.Y(N10898),.A(N10820),.B(N9499));
NAND2X1 NAND2_3275 (.Y(N10899),.A(N10862),.B(N10824));
NAND2X1 NAND2_3276 (.Y(N10902),.A(N10863),.B(N10826));
OR2X1 OR2_3277 (.Y(N10905),.A(N10864),.B(N10765));
OR2X1 OR2_3278 (.Y(N10906),.A(N10865),.B(N10766));
OR2X1 OR2_3279 (.Y(N10907),.A(N10866),.B(N10767));
OR2X1 OR2_3280 (.Y(N10908),.A(N10867),.B(N10768));
NAND2X1 NAND2_3281 (.Y(N10909),.A(N7450),.B(N10872));
NAND2X1 NAND2_3282 (.Y(N10910),.A(N7468),.B(N10874));
NAND2X1 NAND2_3283 (.Y(N10915),.A(N7506),.B(N10882));
NAND2X1 NAND2_3284 (.Y(N10916),.A(N7524),.B(N10884));
NAND2X1 NAND2_3285 (.Y(N10917),.A(N8681),.B(N10886));
NAND2X1 NAND2_3286 (.Y(N10918),.A(N8693),.B(N10888));
NAND2X1 NAND2_3287 (.Y(N10919),.A(N9462),.B(N10890));
NAND2X1 NAND2_3288 (.Y(N10922),.A(N8760),.B(N10895));
NAND2X1 NAND2_3289 (.Y(N10923),.A(N8772),.B(N10897));
NAND2X1 NAND2_3290 (.Y(N10928),.A(N10909),.B(N10873));
NAND2X1 NAND2_3291 (.Y(N10931),.A(N10910),.B(N10875));
INVX1 NOT1_3292 (.Y(N10934),.A(N10876));
NAND2X1 NAND2_3293 (.Y(N10935),.A(N10876),.B(N8634));
INVX1 NOT1_3294 (.Y(N10936),.A(N10879));
NAND2X1 NAND2_3295 (.Y(N10937),.A(N10879),.B(N8639));
NAND2X1 NAND2_3296 (.Y(N10938),.A(N10915),.B(N10883));
NAND2X1 NAND2_3297 (.Y(N10941),.A(N10916),.B(N10885));
NAND2X1 NAND2_3298 (.Y(N10944),.A(N10917),.B(N10887));
NAND2X1 NAND2_3299 (.Y(N10947),.A(N10918),.B(N10889));
NAND2X1 NAND2_3300 (.Y(N10950),.A(N10919),.B(N10891));
INVX1 NOT1_3301 (.Y(N10953),.A(N10892));
NAND2X1 NAND2_3302 (.Y(N10954),.A(N10892),.B(N9476));
NAND2X1 NAND2_3303 (.Y(N10955),.A(N10922),.B(N10896));
NAND2X1 NAND2_3304 (.Y(N10958),.A(N10923),.B(N10898));
INVX1 NOT1_3305 (.Y(N10961),.A(N10899));
NAND2X1 NAND2_3306 (.Y(N10962),.A(N10899),.B(N9506));
INVX1 NOT1_3307 (.Y(N10963),.A(N10902));
NAND2X1 NAND2_3308 (.Y(N10964),.A(N10902),.B(N9515));
NAND2X1 NAND2_3309 (.Y(N10969),.A(N7485),.B(N10934));
NAND2X1 NAND2_3310 (.Y(N10970),.A(N7497),.B(N10936));
NAND2X1 NAND2_3311 (.Y(N10981),.A(N8718),.B(N10953));
NAND2X1 NAND2_3312 (.Y(N10986),.A(N8784),.B(N10961));
NAND2X1 NAND2_3313 (.Y(N10987),.A(N8802),.B(N10963));
INVX1 NOT1_3314 (.Y(N10988),.A(N10928));
NAND2X1 NAND2_3315 (.Y(N10989),.A(N10928),.B(N8617));
INVX1 NOT1_3316 (.Y(N10990),.A(N10931));
NAND2X1 NAND2_3317 (.Y(N10991),.A(N10931),.B(N8626));
NAND2X1 NAND2_3318 (.Y(N10992),.A(N10969),.B(N10935));
NAND2X1 NAND2_3319 (.Y(N10995),.A(N10970),.B(N10937));
INVX1 NOT1_3320 (.Y(N10998),.A(N10938));
NAND2X1 NAND2_3321 (.Y(N10999),.A(N10938),.B(N8646));
INVX1 NOT1_3322 (.Y(N11000),.A(N10941));
NAND2X1 NAND2_3323 (.Y(N11001),.A(N10941),.B(N8655));
INVX1 NOT1_3324 (.Y(N11002),.A(N10944));
NAND2X1 NAND2_3325 (.Y(N11003),.A(N10944),.B(N9456));
INVX1 NOT1_3326 (.Y(N11004),.A(N10947));
NAND2X1 NAND2_3327 (.Y(N11005),.A(N10947),.B(N9461));
INVX1 NOT1_3328 (.Y(N11006),.A(N10950));
NAND2X1 NAND2_3329 (.Y(N11007),.A(N10950),.B(N9465));
NAND2X1 NAND2_3330 (.Y(N11008),.A(N10981),.B(N10954));
INVX1 NOT1_3331 (.Y(N11011),.A(N10955));
NAND2X1 NAND2_3332 (.Y(N11012),.A(N10955),.B(N9495));
INVX1 NOT1_3333 (.Y(N11013),.A(N10958));
NAND2X1 NAND2_3334 (.Y(N11014),.A(N10958),.B(N9500));
NAND2X1 NAND2_3335 (.Y(N11015),.A(N10986),.B(N10962));
NAND2X1 NAND2_3336 (.Y(N11018),.A(N10987),.B(N10964));
NAND2X1 NAND2_3337 (.Y(N11023),.A(N7453),.B(N10988));
NAND2X1 NAND2_3338 (.Y(N11024),.A(N7471),.B(N10990));
NAND2X1 NAND2_3339 (.Y(N11027),.A(N7509),.B(N10998));
NAND2X1 NAND2_3340 (.Y(N11028),.A(N7527),.B(N11000));
NAND2X1 NAND2_3341 (.Y(N11029),.A(N8684),.B(N11002));
NAND2X1 NAND2_3342 (.Y(N11030),.A(N8696),.B(N11004));
NAND2X1 NAND2_3343 (.Y(N11031),.A(N8702),.B(N11006));
NAND2X1 NAND2_3344 (.Y(N11034),.A(N8763),.B(N11011));
NAND2X1 NAND2_3345 (.Y(N11035),.A(N8775),.B(N11013));
INVX1 NOT1_3346 (.Y(N11040),.A(N10992));
NAND2X1 NAND2_3347 (.Y(N11041),.A(N10992),.B(N8294));
INVX1 NOT1_3348 (.Y(N11042),.A(N10995));
NAND2X1 NAND2_3349 (.Y(N11043),.A(N10995),.B(N8295));
NAND2X1 NAND2_3350 (.Y(N11044),.A(N11023),.B(N10989));
NAND2X1 NAND2_3351 (.Y(N11047),.A(N11024),.B(N10991));
NAND2X1 NAND2_3352 (.Y(N11050),.A(N11027),.B(N10999));
NAND2X1 NAND2_3353 (.Y(N11053),.A(N11028),.B(N11001));
NAND2X1 NAND2_3354 (.Y(N11056),.A(N11029),.B(N11003));
NAND2X1 NAND2_3355 (.Y(N11059),.A(N11030),.B(N11005));
NAND2X1 NAND2_3356 (.Y(N11062),.A(N11031),.B(N11007));
INVX1 NOT1_3357 (.Y(N11065),.A(N11008));
NAND2X1 NAND2_3358 (.Y(N11066),.A(N11008),.B(N9477));
NAND2X1 NAND2_3359 (.Y(N11067),.A(N11034),.B(N11012));
NAND2X1 NAND2_3360 (.Y(N11070),.A(N11035),.B(N11014));
INVX1 NOT1_3361 (.Y(N11073),.A(N11015));
NAND2X1 NAND2_3362 (.Y(N11074),.A(N11015),.B(N9507));
INVX1 NOT1_3363 (.Y(N11075),.A(N11018));
NAND2X1 NAND2_3364 (.Y(N11076),.A(N11018),.B(N9516));
NAND2X1 NAND2_3365 (.Y(N11077),.A(N7488),.B(N11040));
NAND2X1 NAND2_3366 (.Y(N11078),.A(N7500),.B(N11042));
NAND2X1 NAND2_3367 (.Y(N11095),.A(N8721),.B(N11065));
NAND2X1 NAND2_3368 (.Y(N11098),.A(N8787),.B(N11073));
NAND2X1 NAND2_3369 (.Y(N11099),.A(N8805),.B(N11075));
NAND2X1 NAND2_3370 (.Y(N11100),.A(N11077),.B(N11041));
NAND2X1 NAND2_3371 (.Y(N11103),.A(N11078),.B(N11043));
INVX1 NOT1_3372 (.Y(N11106),.A(N11056));
NAND2X1 NAND2_3373 (.Y(N11107),.A(N11056),.B(N9319));
INVX1 NOT1_3374 (.Y(N11108),.A(N11059));
NAND2X1 NAND2_3375 (.Y(N11109),.A(N11059),.B(N9320));
INVX1 NOT1_3376 (.Y(N11110),.A(N11067));
NAND2X1 NAND2_3377 (.Y(N11111),.A(N11067),.B(N9381));
INVX1 NOT1_3378 (.Y(N11112),.A(N11070));
NAND2X1 NAND2_3379 (.Y(N11113),.A(N11070),.B(N9382));
INVX1 NOT1_3380 (.Y(N11114),.A(N11044));
NAND2X1 NAND2_3381 (.Y(N11115),.A(N11044),.B(N8618));
INVX1 NOT1_3382 (.Y(N11116),.A(N11047));
NAND2X1 NAND2_3383 (.Y(N11117),.A(N11047),.B(N8619));
INVX1 NOT1_3384 (.Y(N11118),.A(N11050));
NAND2X1 NAND2_3385 (.Y(N11119),.A(N11050),.B(N8647));
INVX1 NOT1_3386 (.Y(N11120),.A(N11053));
NAND2X1 NAND2_3387 (.Y(N11121),.A(N11053),.B(N8648));
INVX1 NOT1_3388 (.Y(N11122),.A(N11062));
NAND2X1 NAND2_3389 (.Y(N11123),.A(N11062),.B(N9466));
NAND2X1 NAND2_3390 (.Y(N11124),.A(N11095),.B(N11066));
NAND2X1 NAND2_3391 (.Y(N11127),.A(N11098),.B(N11074));
NAND2X1 NAND2_3392 (.Y(N11130),.A(N11099),.B(N11076));
NAND2X1 NAND2_3393 (.Y(N11137),.A(N8687),.B(N11106));
NAND2X1 NAND2_3394 (.Y(N11138),.A(N8699),.B(N11108));
NAND2X1 NAND2_3395 (.Y(N11139),.A(N8766),.B(N11110));
NAND2X1 NAND2_3396 (.Y(N11140),.A(N8778),.B(N11112));
NAND2X1 NAND2_3397 (.Y(N11141),.A(N7456),.B(N11114));
NAND2X1 NAND2_3398 (.Y(N11142),.A(N7474),.B(N11116));
NAND2X1 NAND2_3399 (.Y(N11143),.A(N7512),.B(N11118));
NAND2X1 NAND2_3400 (.Y(N11144),.A(N7530),.B(N11120));
NAND2X1 NAND2_3401 (.Y(N11145),.A(N8705),.B(N11122));
AND2X1 AND_tmp818 (.Y(ttmp818),.A(N8871),.B(N10283));
AND2X1 AND_tmp819 (.Y(N11152),.A(N11103),.B(ttmp818));
AND2X1 AND_tmp820 (.Y(ttmp820),.A(N7655),.B(N10283));
AND2X1 AND_tmp821 (.Y(N11153),.A(N11100),.B(ttmp820));
AND2X1 AND_tmp822 (.Y(ttmp822),.A(N9551),.B(N10119));
AND2X1 AND_tmp823 (.Y(N11154),.A(N11103),.B(ttmp822));
AND2X1 AND_tmp824 (.Y(ttmp824),.A(N9917),.B(N10119));
AND2X1 AND_tmp825 (.Y(N11155),.A(N11100),.B(ttmp824));
NAND2X1 NAND2_3406 (.Y(N11156),.A(N11137),.B(N11107));
NAND2X1 NAND2_3407 (.Y(N11159),.A(N11138),.B(N11109));
NAND2X1 NAND2_3408 (.Y(N11162),.A(N11139),.B(N11111));
NAND2X1 NAND2_3409 (.Y(N11165),.A(N11140),.B(N11113));
NAND2X1 NAND2_3410 (.Y(N11168),.A(N11141),.B(N11115));
NAND2X1 NAND2_3411 (.Y(N11171),.A(N11142),.B(N11117));
NAND2X1 NAND2_3412 (.Y(N11174),.A(N11143),.B(N11119));
NAND2X1 NAND2_3413 (.Y(N11177),.A(N11144),.B(N11121));
NAND2X1 NAND2_3414 (.Y(N11180),.A(N11145),.B(N11123));
INVX1 NOT1_3415 (.Y(N11183),.A(N11124));
NAND2X1 NAND2_3416 (.Y(N11184),.A(N11124),.B(N9468));
INVX1 NOT1_3417 (.Y(N11185),.A(N11127));
NAND2X1 NAND2_3418 (.Y(N11186),.A(N11127),.B(N9508));
INVX1 NOT1_3419 (.Y(N11187),.A(N11130));
NAND2X1 NAND2_3420 (.Y(N11188),.A(N11130),.B(N9509));
OR2X1 OR_tmp826 (.Y(ttmp826),.A(N11154),.B(N11155));
OR2X1 OR_tmp827 (.Y(ttmp827),.A(N11152),.B(ttmp826));
OR2X1 OR_tmp828 (.Y(N11205),.A(N11153),.B(ttmp827));
NAND2X1 NAND2_3422 (.Y(N11210),.A(N8724),.B(N11183));
NAND2X1 NAND2_3423 (.Y(N11211),.A(N8790),.B(N11185));
NAND2X1 NAND2_3424 (.Y(N11212),.A(N8808),.B(N11187));
INVX1 NOT1_3425 (.Y(N11213),.A(N11168));
NAND2X1 NAND2_3426 (.Y(N11214),.A(N11168),.B(N8260));
INVX1 NOT1_3427 (.Y(N11215),.A(N11171));
NAND2X1 NAND2_3428 (.Y(N11216),.A(N11171),.B(N8261));
INVX1 NOT1_3429 (.Y(N11217),.A(N11174));
NAND2X1 NAND2_3430 (.Y(N11218),.A(N11174),.B(N8296));
INVX1 NOT1_3431 (.Y(N11219),.A(N11177));
NAND2X1 NAND2_3432 (.Y(N11220),.A(N11177),.B(N8297));
AND2X1 AND_tmp829 (.Y(ttmp829),.A(N9575),.B(N1218));
AND2X1 AND_tmp830 (.Y(N11222),.A(N11159),.B(ttmp829));
AND2X1 AND_tmp831 (.Y(ttmp831),.A(N8927),.B(N1218));
AND2X1 AND_tmp832 (.Y(N11223),.A(N11156),.B(ttmp831));
AND2X1 AND_tmp833 (.Y(ttmp833),.A(N9935),.B(N750));
AND2X1 AND_tmp834 (.Y(N11224),.A(N11159),.B(ttmp833));
AND2X1 AND_tmp835 (.Y(ttmp835),.A(N10132),.B(N750));
AND2X1 AND_tmp836 (.Y(N11225),.A(N11156),.B(ttmp835));
AND2X1 AND_tmp837 (.Y(ttmp837),.A(N9608),.B(N10497));
AND2X1 AND_tmp838 (.Y(N11226),.A(N11165),.B(ttmp837));
AND2X1 AND_tmp839 (.Y(ttmp839),.A(N9001),.B(N10497));
AND2X1 AND_tmp840 (.Y(N11227),.A(N11162),.B(ttmp839));
AND2X1 AND_tmp841 (.Y(ttmp841),.A(N9949),.B(N10301));
AND2X1 AND_tmp842 (.Y(N11228),.A(N11165),.B(ttmp841));
AND2X1 AND_tmp843 (.Y(ttmp843),.A(N10160),.B(N10301));
AND2X1 AND_tmp844 (.Y(N11229),.A(N11162),.B(ttmp843));
INVX1 NOT1_3441 (.Y(N11231),.A(N11180));
NAND2X1 NAND2_3442 (.Y(N11232),.A(N11180),.B(N9467));
NAND2X1 NAND2_3443 (.Y(N11233),.A(N11210),.B(N11184));
NAND2X1 NAND2_3444 (.Y(N11236),.A(N11211),.B(N11186));
NAND2X1 NAND2_3445 (.Y(N11239),.A(N11212),.B(N11188));
NAND2X1 NAND2_3446 (.Y(N11242),.A(N7459),.B(N11213));
NAND2X1 NAND2_3447 (.Y(N11243),.A(N7462),.B(N11215));
NAND2X1 NAND2_3448 (.Y(N11244),.A(N7515),.B(N11217));
NAND2X1 NAND2_3449 (.Y(N11245),.A(N7518),.B(N11219));
INVX1 NOT1_3450 (.Y(N11246),.A(N11205));
NAND2X1 NAND2_3451 (.Y(N11250),.A(N8708),.B(N11231));
OR2X1 OR_tmp845 (.Y(ttmp845),.A(N11224),.B(N11225));
OR2X1 OR_tmp846 (.Y(ttmp846),.A(N11222),.B(ttmp845));
OR2X1 OR_tmp847 (.Y(N11252),.A(N11223),.B(ttmp846));
OR2X1 OR_tmp848 (.Y(ttmp848),.A(N11228),.B(N11229));
OR2X1 OR_tmp849 (.Y(ttmp849),.A(N11226),.B(ttmp848));
OR2X1 OR_tmp850 (.Y(N11257),.A(N11227),.B(ttmp849));
NAND2X1 NAND2_3454 (.Y(N11260),.A(N11242),.B(N11214));
NAND2X1 NAND2_3455 (.Y(N11261),.A(N11243),.B(N11216));
NAND2X1 NAND2_3456 (.Y(N11262),.A(N11244),.B(N11218));
NAND2X1 NAND2_3457 (.Y(N11263),.A(N11245),.B(N11220));
INVX1 NOT1_3458 (.Y(N11264),.A(N11233));
NAND2X1 NAND2_3459 (.Y(N11265),.A(N11233),.B(N9322));
INVX1 NOT1_3460 (.Y(N11267),.A(N11236));
NAND2X1 NAND2_3461 (.Y(N11268),.A(N11236),.B(N9383));
INVX1 NOT1_3462 (.Y(N11269),.A(N11239));
NAND2X1 NAND2_3463 (.Y(N11270),.A(N11239),.B(N9384));
NAND2X1 NAND2_3464 (.Y(N11272),.A(N11250),.B(N11232));
INVX1 NOT1_3465 (.Y(N11277),.A(N11261));
AND2X1 AND2_3466 (.Y(N11278),.A(N10273),.B(N11260));
INVX1 NOT1_3467 (.Y(N11279),.A(N11263));
AND2X1 AND2_3468 (.Y(N11280),.A(N10119),.B(N11262));
NAND2X1 NAND2_3469 (.Y(N11282),.A(N8714),.B(N11264));
INVX1 NOT1_3470 (.Y(N11283),.A(N11252));
NAND2X1 NAND2_3471 (.Y(N11284),.A(N8793),.B(N11267));
NAND2X1 NAND2_3472 (.Y(N11285),.A(N8796),.B(N11269));
INVX1 NOT1_3473 (.Y(N11286),.A(N11257));
AND2X1 AND2_3474 (.Y(N11288),.A(N11277),.B(N10479));
AND2X1 AND2_3475 (.Y(N11289),.A(N11279),.B(N10283));
INVX1 NOT1_3476 (.Y(N11290),.A(N11272));
NAND2X1 NAND2_3477 (.Y(N11291),.A(N11272),.B(N9321));
NAND2X1 NAND2_3478 (.Y(N11292),.A(N11282),.B(N11265));
NAND2X1 NAND2_3479 (.Y(N11293),.A(N11284),.B(N11268));
NAND2X1 NAND2_3480 (.Y(N11294),.A(N11285),.B(N11270));
NAND2X1 NAND2_3481 (.Y(N11295),.A(N8711),.B(N11290));
INVX1 NOT1_3482 (.Y(N11296),.A(N11292));
INVX1 NOT1_3483 (.Y(N11297),.A(N11294));
AND2X1 AND2_3484 (.Y(N11298),.A(N10301),.B(N11293));
OR2X1 OR2_3485 (.Y(N11299),.A(N11288),.B(N11278));
OR2X1 OR2_3486 (.Y(N11302),.A(N11289),.B(N11280));
NAND2X1 NAND2_3487 (.Y(N11307),.A(N11295),.B(N11291));
AND2X1 AND2_3488 (.Y(N11308),.A(N11296),.B(N1218));
AND2X1 AND2_3489 (.Y(N11309),.A(N11297),.B(N10497));
NAND2X1 NAND2_3490 (.Y(N11312),.A(N11302),.B(N11246));
NAND2X1 NAND2_3491 (.Y(N11313),.A(N11299),.B(N10836));
INVX1 NOT1_3492 (.Y(N11314),.A(N11299));
INVX1 NOT1_3493 (.Y(N11315),.A(N11302));
AND2X1 AND2_3494 (.Y(N11316),.A(N750),.B(N11307));
OR2X1 OR2_3495 (.Y(N11317),.A(N11309),.B(N11298));
NAND2X1 NAND2_3496 (.Y(N11320),.A(N11205),.B(N11315));
NAND2X1 NAND2_3497 (.Y(N11321),.A(N10739),.B(N11314));
OR2X1 OR2_3498 (.Y(N11323),.A(N11308),.B(N11316));
NAND2X1 NAND2_3499 (.Y(N11327),.A(N11312),.B(N11320));
NAND2X1 NAND2_3500 (.Y(N11328),.A(N11313),.B(N11321));
NAND2X1 NAND2_3501 (.Y(N11329),.A(N11317),.B(N11286));
INVX1 NOT1_3502 (.Y(N11331),.A(N11317));
INVX1 NOT1_3503 (.Y(N11333),.A(N11327));
INVX1 NOT1_3504 (.Y(N11334),.A(N11328));
NAND2X1 NAND2_3505 (.Y(N11335),.A(N11257),.B(N11331));
NAND2X1 NAND2_3506 (.Y(N11336),.A(N11323),.B(N11283));
INVX1 NOT1_3507 (.Y(N11337),.A(N11323));
NAND2X1 NAND2_3508 (.Y(N11338),.A(N11329),.B(N11335));
NAND2X1 NAND2_3509 (.Y(N11339),.A(N11252),.B(N11337));
INVX1 NOT1_3510 (.Y(N11340),.A(N11338));
NAND2X1 NAND2_3511 (.Y(N11341),.A(N11336),.B(N11339));
INVX1 NOT1_3512 (.Y(N11342),.A(N11341));
BUFX1 BUFF1_3513 (.Y(N241_O),.A(N241_I));
endmodule