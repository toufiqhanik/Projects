module c17 (N1,N2,N3,N6,N7,N22,N23,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9);
input N1,N2,N3,N6,N7,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9;
output N22,N23;
wire N10,N11,N16,N19,N7enc,N3enc,N19enc,N16enc,N22enc,xorgate0,xorgate1,xorgate2,xorgate3,xorgate4,compare0,compare1,compare2,compare3,compare4,andgate0,andgate1,andgate2,andgate3,orgate0,orgate1,orgate2,orgate3,andgate4,N22_sar,N23_sar;
NAND2X1 NAND2_1 (.Y(N10),.A(N1),.B(N3enc));
NAND2X1 NAND2_2 (.Y(N11),.A(N3enc),.B(N6));
NAND2X1 NAND2_3 (.Y(N16),.A(N2),.B(N11));
NAND2X1 NAND2_4 (.Y(N19),.A(N11),.B(N7enc));
NAND2X1 NAND2_5 (.Y(N22enc),.A(N10),.B(N16enc));
NAND2X1 NAND2_6 (.Y(N23_sar),.A(N16enc),.B(N19enc));
XOR2X1 XOR2_N7 (.Y(N7enc),.A(N7),.B(keyinput0));
XNOR2X1 XNOR2_N3 (.Y(N3enc),.A(N3),.B(keyinput1));
XOR2X1 XOR2_N19 (.Y(N19enc),.A(N19),.B(keyinput2));
XNOR2X1 XNOR2_N16 (.Y(N16enc),.A(N16),.B(keyinput3));
XNOR2X1 XNOR2_N22 (.Y(N22_sar),.A(N22enc),.B(keyinput4));
XOR2X1 xorgate_0 (.Y(xorgate0),.A(keyinput0),.B(keyinput5));
XOR2X1 xorgate_1 (.Y(xorgate1),.A(keyinput1),.B(keyinput6));
XOR2X1 xorgate_2 (.Y(xorgate2),.A(keyinput2),.B(keyinput7));
XOR2X1 xorgate_3 (.Y(xorgate3),.A(keyinput3),.B(keyinput8));
XOR2X1 xorgate_4 (.Y(xorgate4),.A(keyinput4),.B(keyinput9));
XNOR2X1 compare_0 (.Y(compare0),.A(xorgate0),.B(N1));
XNOR2X1 compare_1 (.Y(compare1),.A(xorgate1),.B(N2));
XNOR2X1 compare_2 (.Y(compare2),.A(xorgate2),.B(N3));
XNOR2X1 compare_3 (.Y(compare3),.A(xorgate3),.B(N6));
XNOR2X1 compare_4 (.Y(compare4),.A(xorgate4),.B(N7));
AND2X1 andgate_0 (.Y(andgate0),.A(compare0),.B(compare1));
AND2X1 andgate_1 (.Y(andgate1),.A(compare2),.B(compare3));
AND2X1 andgate_2 (.Y(andgate2),.A(compare4),.B(andgate0));
AND2X1 andgate_3 (.Y(andgate3),.A(andgate1),.B(andgate2));
OR2X1 orgate_0 (.Y(orgate0),.A(keyinput5),.B(keyinput6));
OR2X1 orgate_1 (.Y(orgate1),.A(keyinput7),.B(keyinput8));
OR2X1 orgate_2 (.Y(orgate2),.A(keyinput9),.B(orgate0));
OR2X1 orgate_3 (.Y(orgate3),.A(orgate1),.B(orgate2));
AND2X1 andgate_4 (.Y(andgate4),.A(orgate3),.B(andgate3));
XOR2X1 XOR_out0 (.Y(N22),.A(N22_sar),.B(andgate4));
XOR2X1 XOR_out1 (.Y(N23),.A(N23_sar),.B(andgate4));
endmodule