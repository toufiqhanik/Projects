module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755);
input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,N137;
output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755;
wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723;
XOR2X1 XOR2_1 (.Y(N250),.A(N1),.B(N5));
XOR2X1 XOR2_2 (.Y(N251),.A(N9),.B(N13));
XOR2X1 XOR2_3 (.Y(N252),.A(N17),.B(N21));
XOR2X1 XOR2_4 (.Y(N253),.A(N25),.B(N29));
XOR2X1 XOR2_5 (.Y(N254),.A(N33),.B(N37));
XOR2X1 XOR2_6 (.Y(N255),.A(N41),.B(N45));
XOR2X1 XOR2_7 (.Y(N256),.A(N49),.B(N53));
XOR2X1 XOR2_8 (.Y(N257),.A(N57),.B(N61));
XOR2X1 XOR2_9 (.Y(N258),.A(N65),.B(N69));
XOR2X1 XOR2_10 (.Y(N259),.A(N73),.B(N77));
XOR2X1 XOR2_11 (.Y(N260),.A(N81),.B(N85));
XOR2X1 XOR2_12 (.Y(N261),.A(N89),.B(N93));
XOR2X1 XOR2_13 (.Y(N262),.A(N97),.B(N101));
XOR2X1 XOR2_14 (.Y(N263),.A(N105),.B(N109));
XOR2X1 XOR2_15 (.Y(N264),.A(N113),.B(N117));
XOR2X1 XOR2_16 (.Y(N265),.A(N121),.B(N125));
AND2X1 AND2_17 (.Y(N266),.A(N129),.B(N137));
AND2X1 AND2_18 (.Y(N267),.A(N130),.B(N137));
AND2X1 AND2_19 (.Y(N268),.A(N131),.B(N137));
AND2X1 AND2_20 (.Y(N269),.A(N132),.B(N137));
AND2X1 AND2_21 (.Y(N270),.A(N133),.B(N137));
AND2X1 AND2_22 (.Y(N271),.A(N134),.B(N137));
AND2X1 AND2_23 (.Y(N272),.A(N135),.B(N137));
AND2X1 AND2_24 (.Y(N273),.A(N136),.B(N137));
XOR2X1 XOR2_25 (.Y(N274),.A(N1),.B(N17));
XOR2X1 XOR2_26 (.Y(N275),.A(N33),.B(N49));
XOR2X1 XOR2_27 (.Y(N276),.A(N5),.B(N21));
XOR2X1 XOR2_28 (.Y(N277),.A(N37),.B(N53));
XOR2X1 XOR2_29 (.Y(N278),.A(N9),.B(N25));
XOR2X1 XOR2_30 (.Y(N279),.A(N41),.B(N57));
XOR2X1 XOR2_31 (.Y(N280),.A(N13),.B(N29));
XOR2X1 XOR2_32 (.Y(N281),.A(N45),.B(N61));
XOR2X1 XOR2_33 (.Y(N282),.A(N65),.B(N81));
XOR2X1 XOR2_34 (.Y(N283),.A(N97),.B(N113));
XOR2X1 XOR2_35 (.Y(N284),.A(N69),.B(N85));
XOR2X1 XOR2_36 (.Y(N285),.A(N101),.B(N117));
XOR2X1 XOR2_37 (.Y(N286),.A(N73),.B(N89));
XOR2X1 XOR2_38 (.Y(N287),.A(N105),.B(N121));
XOR2X1 XOR2_39 (.Y(N288),.A(N77),.B(N93));
XOR2X1 XOR2_40 (.Y(N289),.A(N109),.B(N125));
XOR2X1 XOR2_41 (.Y(N290),.A(N250),.B(N251));
XOR2X1 XOR2_42 (.Y(N293),.A(N252),.B(N253));
XOR2X1 XOR2_43 (.Y(N296),.A(N254),.B(N255));
XOR2X1 XOR2_44 (.Y(N299),.A(N256),.B(N257));
XOR2X1 XOR2_45 (.Y(N302),.A(N258),.B(N259));
XOR2X1 XOR2_46 (.Y(N305),.A(N260),.B(N261));
XOR2X1 XOR2_47 (.Y(N308),.A(N262),.B(N263));
XOR2X1 XOR2_48 (.Y(N311),.A(N264),.B(N265));
XOR2X1 XOR2_49 (.Y(N314),.A(N274),.B(N275));
XOR2X1 XOR2_50 (.Y(N315),.A(N276),.B(N277));
XOR2X1 XOR2_51 (.Y(N316),.A(N278),.B(N279));
XOR2X1 XOR2_52 (.Y(N317),.A(N280),.B(N281));
XOR2X1 XOR2_53 (.Y(N318),.A(N282),.B(N283));
XOR2X1 XOR2_54 (.Y(N319),.A(N284),.B(N285));
XOR2X1 XOR2_55 (.Y(N320),.A(N286),.B(N287));
XOR2X1 XOR2_56 (.Y(N321),.A(N288),.B(N289));
XOR2X1 XOR2_57 (.Y(N338),.A(N290),.B(N293));
XOR2X1 XOR2_58 (.Y(N339),.A(N296),.B(N299));
XOR2X1 XOR2_59 (.Y(N340),.A(N290),.B(N296));
XOR2X1 XOR2_60 (.Y(N341),.A(N293),.B(N299));
XOR2X1 XOR2_61 (.Y(N342),.A(N302),.B(N305));
XOR2X1 XOR2_62 (.Y(N343),.A(N308),.B(N311));
XOR2X1 XOR2_63 (.Y(N344),.A(N302),.B(N308));
XOR2X1 XOR2_64 (.Y(N345),.A(N305),.B(N311));
XOR2X1 XOR2_65 (.Y(N346),.A(N266),.B(N342));
XOR2X1 XOR2_66 (.Y(N347),.A(N267),.B(N343));
XOR2X1 XOR2_67 (.Y(N348),.A(N268),.B(N344));
XOR2X1 XOR2_68 (.Y(N349),.A(N269),.B(N345));
XOR2X1 XOR2_69 (.Y(N350),.A(N270),.B(N338));
XOR2X1 XOR2_70 (.Y(N351),.A(N271),.B(N339));
XOR2X1 XOR2_71 (.Y(N352),.A(N272),.B(N340));
XOR2X1 XOR2_72 (.Y(N353),.A(N273),.B(N341));
XOR2X1 XOR2_73 (.Y(N354),.A(N314),.B(N346));
XOR2X1 XOR2_74 (.Y(N367),.A(N315),.B(N347));
XOR2X1 XOR2_75 (.Y(N380),.A(N316),.B(N348));
XOR2X1 XOR2_76 (.Y(N393),.A(N317),.B(N349));
XOR2X1 XOR2_77 (.Y(N406),.A(N318),.B(N350));
XOR2X1 XOR2_78 (.Y(N419),.A(N319),.B(N351));
XOR2X1 XOR2_79 (.Y(N432),.A(N320),.B(N352));
XOR2X1 XOR2_80 (.Y(N445),.A(N321),.B(N353));
INVX1 NOT1_81 (.Y(N554),.A(N354));
INVX1 NOT1_82 (.Y(N555),.A(N367));
INVX1 NOT1_83 (.Y(N556),.A(N380));
INVX1 NOT1_84 (.Y(N557),.A(N354));
INVX1 NOT1_85 (.Y(N558),.A(N367));
INVX1 NOT1_86 (.Y(N559),.A(N393));
INVX1 NOT1_87 (.Y(N560),.A(N354));
INVX1 NOT1_88 (.Y(N561),.A(N380));
INVX1 NOT1_89 (.Y(N562),.A(N393));
INVX1 NOT1_90 (.Y(N563),.A(N367));
INVX1 NOT1_91 (.Y(N564),.A(N380));
INVX1 NOT1_92 (.Y(N565),.A(N393));
INVX1 NOT1_93 (.Y(N566),.A(N419));
INVX1 NOT1_94 (.Y(N567),.A(N445));
INVX1 NOT1_95 (.Y(N568),.A(N419));
INVX1 NOT1_96 (.Y(N569),.A(N432));
INVX1 NOT1_97 (.Y(N570),.A(N406));
INVX1 NOT1_98 (.Y(N571),.A(N445));
INVX1 NOT1_99 (.Y(N572),.A(N406));
INVX1 NOT1_100 (.Y(N573),.A(N432));
INVX1 NOT1_101 (.Y(N574),.A(N406));
INVX1 NOT1_102 (.Y(N575),.A(N419));
INVX1 NOT1_103 (.Y(N576),.A(N432));
INVX1 NOT1_104 (.Y(N577),.A(N406));
INVX1 NOT1_105 (.Y(N578),.A(N419));
INVX1 NOT1_106 (.Y(N579),.A(N445));
INVX1 NOT1_107 (.Y(N580),.A(N406));
INVX1 NOT1_108 (.Y(N581),.A(N432));
INVX1 NOT1_109 (.Y(N582),.A(N445));
INVX1 NOT1_110 (.Y(N583),.A(N419));
INVX1 NOT1_111 (.Y(N584),.A(N432));
INVX1 NOT1_112 (.Y(N585),.A(N445));
INVX1 NOT1_113 (.Y(N586),.A(N367));
INVX1 NOT1_114 (.Y(N587),.A(N393));
INVX1 NOT1_115 (.Y(N588),.A(N367));
INVX1 NOT1_116 (.Y(N589),.A(N380));
INVX1 NOT1_117 (.Y(N590),.A(N354));
INVX1 NOT1_118 (.Y(N591),.A(N393));
INVX1 NOT1_119 (.Y(N592),.A(N354));
INVX1 NOT1_120 (.Y(N593),.A(N380));
AND2X1 AND_tmp1 (.Y(ttmp1),.A(N556),.B(N393));
AND2X1 AND_tmp2 (.Y(ttmp2),.A(N554),.B(ttmp1));
AND2X1 AND_tmp3 (.Y(N594),.A(N555),.B(ttmp2));
AND2X1 AND_tmp4 (.Y(ttmp4),.A(N380),.B(N559));
AND2X1 AND_tmp5 (.Y(ttmp5),.A(N557),.B(ttmp4));
AND2X1 AND_tmp6 (.Y(N595),.A(N558),.B(ttmp5));
AND2X1 AND_tmp7 (.Y(ttmp7),.A(N561),.B(N562));
AND2X1 AND_tmp8 (.Y(ttmp8),.A(N560),.B(ttmp7));
AND2X1 AND_tmp9 (.Y(N596),.A(N367),.B(ttmp8));
AND2X1 AND_tmp10 (.Y(ttmp10),.A(N564),.B(N565));
AND2X1 AND_tmp11 (.Y(ttmp11),.A(N354),.B(ttmp10));
AND2X1 AND_tmp12 (.Y(N597),.A(N563),.B(ttmp11));
AND2X1 AND_tmp13 (.Y(ttmp13),.A(N576),.B(N445));
AND2X1 AND_tmp14 (.Y(ttmp14),.A(N574),.B(ttmp13));
AND2X1 AND_tmp15 (.Y(N598),.A(N575),.B(ttmp14));
AND2X1 AND_tmp16 (.Y(ttmp16),.A(N432),.B(N579));
AND2X1 AND_tmp17 (.Y(ttmp17),.A(N577),.B(ttmp16));
AND2X1 AND_tmp18 (.Y(N599),.A(N578),.B(ttmp17));
AND2X1 AND_tmp19 (.Y(ttmp19),.A(N581),.B(N582));
AND2X1 AND_tmp20 (.Y(ttmp20),.A(N580),.B(ttmp19));
AND2X1 AND_tmp21 (.Y(N600),.A(N419),.B(ttmp20));
AND2X1 AND_tmp22 (.Y(ttmp22),.A(N584),.B(N585));
AND2X1 AND_tmp23 (.Y(ttmp23),.A(N406),.B(ttmp22));
AND2X1 AND_tmp24 (.Y(N601),.A(N583),.B(ttmp23));
OR2X1 OR_tmp25 (.Y(ttmp25),.A(N596),.B(N597));
OR2X1 OR_tmp26 (.Y(ttmp26),.A(N594),.B(ttmp25));
OR2X1 OR_tmp27 (.Y(N602),.A(N595),.B(ttmp26));
OR2X1 OR_tmp28 (.Y(ttmp28),.A(N600),.B(N601));
OR2X1 OR_tmp29 (.Y(ttmp29),.A(N598),.B(ttmp28));
OR2X1 OR_tmp30 (.Y(N607),.A(N599),.B(ttmp29));
AND2X1 AND_tmp31 (.Y(ttmp31),.A(N567),.B(N602));
AND2X1 AND_tmp32 (.Y(ttmp32),.A(N406),.B(ttmp31));
AND2X1 AND_tmp33 (.Y(ttmp33),.A(N566),.B(ttmp32));
AND2X1 AND_tmp34 (.Y(N620),.A(N432),.B(ttmp33));
AND2X1 AND_tmp35 (.Y(ttmp35),.A(N445),.B(N602));
AND2X1 AND_tmp36 (.Y(ttmp36),.A(N406),.B(ttmp35));
AND2X1 AND_tmp37 (.Y(ttmp37),.A(N568),.B(ttmp36));
AND2X1 AND_tmp38 (.Y(N625),.A(N569),.B(ttmp37));
AND2X1 AND_tmp39 (.Y(ttmp39),.A(N571),.B(N602));
AND2X1 AND_tmp40 (.Y(ttmp40),.A(N570),.B(ttmp39));
AND2X1 AND_tmp41 (.Y(ttmp41),.A(N419),.B(ttmp40));
AND2X1 AND_tmp42 (.Y(N630),.A(N432),.B(ttmp41));
AND2X1 AND_tmp43 (.Y(ttmp43),.A(N445),.B(N602));
AND2X1 AND_tmp44 (.Y(ttmp44),.A(N572),.B(ttmp43));
AND2X1 AND_tmp45 (.Y(ttmp45),.A(N419),.B(ttmp44));
AND2X1 AND_tmp46 (.Y(N635),.A(N573),.B(ttmp45));
AND2X1 AND_tmp47 (.Y(ttmp47),.A(N587),.B(N607));
AND2X1 AND_tmp48 (.Y(ttmp48),.A(N354),.B(ttmp47));
AND2X1 AND_tmp49 (.Y(ttmp49),.A(N586),.B(ttmp48));
AND2X1 AND_tmp50 (.Y(N640),.A(N380),.B(ttmp49));
AND2X1 AND_tmp51 (.Y(ttmp51),.A(N393),.B(N607));
AND2X1 AND_tmp52 (.Y(ttmp52),.A(N354),.B(ttmp51));
AND2X1 AND_tmp53 (.Y(ttmp53),.A(N588),.B(ttmp52));
AND2X1 AND_tmp54 (.Y(N645),.A(N589),.B(ttmp53));
AND2X1 AND_tmp55 (.Y(ttmp55),.A(N591),.B(N607));
AND2X1 AND_tmp56 (.Y(ttmp56),.A(N590),.B(ttmp55));
AND2X1 AND_tmp57 (.Y(ttmp57),.A(N367),.B(ttmp56));
AND2X1 AND_tmp58 (.Y(N650),.A(N380),.B(ttmp57));
AND2X1 AND_tmp59 (.Y(ttmp59),.A(N393),.B(N607));
AND2X1 AND_tmp60 (.Y(ttmp60),.A(N592),.B(ttmp59));
AND2X1 AND_tmp61 (.Y(ttmp61),.A(N367),.B(ttmp60));
AND2X1 AND_tmp62 (.Y(N655),.A(N593),.B(ttmp61));
AND2X1 AND2_139 (.Y(N692),.A(N354),.B(N620));
AND2X1 AND2_140 (.Y(N693),.A(N367),.B(N620));
AND2X1 AND2_141 (.Y(N694),.A(N380),.B(N620));
AND2X1 AND2_142 (.Y(N695),.A(N393),.B(N620));
AND2X1 AND2_143 (.Y(N696),.A(N354),.B(N625));
AND2X1 AND2_144 (.Y(N697),.A(N367),.B(N625));
AND2X1 AND2_145 (.Y(N698),.A(N380),.B(N625));
AND2X1 AND2_146 (.Y(N699),.A(N393),.B(N625));
AND2X1 AND2_147 (.Y(N700),.A(N354),.B(N630));
AND2X1 AND2_148 (.Y(N701),.A(N367),.B(N630));
AND2X1 AND2_149 (.Y(N702),.A(N380),.B(N630));
AND2X1 AND2_150 (.Y(N703),.A(N393),.B(N630));
AND2X1 AND2_151 (.Y(N704),.A(N354),.B(N635));
AND2X1 AND2_152 (.Y(N705),.A(N367),.B(N635));
AND2X1 AND2_153 (.Y(N706),.A(N380),.B(N635));
AND2X1 AND2_154 (.Y(N707),.A(N393),.B(N635));
AND2X1 AND2_155 (.Y(N708),.A(N406),.B(N640));
AND2X1 AND2_156 (.Y(N709),.A(N419),.B(N640));
AND2X1 AND2_157 (.Y(N710),.A(N432),.B(N640));
AND2X1 AND2_158 (.Y(N711),.A(N445),.B(N640));
AND2X1 AND2_159 (.Y(N712),.A(N406),.B(N645));
AND2X1 AND2_160 (.Y(N713),.A(N419),.B(N645));
AND2X1 AND2_161 (.Y(N714),.A(N432),.B(N645));
AND2X1 AND2_162 (.Y(N715),.A(N445),.B(N645));
AND2X1 AND2_163 (.Y(N716),.A(N406),.B(N650));
AND2X1 AND2_164 (.Y(N717),.A(N419),.B(N650));
AND2X1 AND2_165 (.Y(N718),.A(N432),.B(N650));
AND2X1 AND2_166 (.Y(N719),.A(N445),.B(N650));
AND2X1 AND2_167 (.Y(N720),.A(N406),.B(N655));
AND2X1 AND2_168 (.Y(N721),.A(N419),.B(N655));
AND2X1 AND2_169 (.Y(N722),.A(N432),.B(N655));
AND2X1 AND2_170 (.Y(N723),.A(N445),.B(N655));
XOR2X1 XOR2_171 (.Y(N724),.A(N1),.B(N692));
XOR2X1 XOR2_172 (.Y(N725),.A(N5),.B(N693));
XOR2X1 XOR2_173 (.Y(N726),.A(N9),.B(N694));
XOR2X1 XOR2_174 (.Y(N727),.A(N13),.B(N695));
XOR2X1 XOR2_175 (.Y(N728),.A(N17),.B(N696));
XOR2X1 XOR2_176 (.Y(N729),.A(N21),.B(N697));
XOR2X1 XOR2_177 (.Y(N730),.A(N25),.B(N698));
XOR2X1 XOR2_178 (.Y(N731),.A(N29),.B(N699));
XOR2X1 XOR2_179 (.Y(N732),.A(N33),.B(N700));
XOR2X1 XOR2_180 (.Y(N733),.A(N37),.B(N701));
XOR2X1 XOR2_181 (.Y(N734),.A(N41),.B(N702));
XOR2X1 XOR2_182 (.Y(N735),.A(N45),.B(N703));
XOR2X1 XOR2_183 (.Y(N736),.A(N49),.B(N704));
XOR2X1 XOR2_184 (.Y(N737),.A(N53),.B(N705));
XOR2X1 XOR2_185 (.Y(N738),.A(N57),.B(N706));
XOR2X1 XOR2_186 (.Y(N739),.A(N61),.B(N707));
XOR2X1 XOR2_187 (.Y(N740),.A(N65),.B(N708));
XOR2X1 XOR2_188 (.Y(N741),.A(N69),.B(N709));
XOR2X1 XOR2_189 (.Y(N742),.A(N73),.B(N710));
XOR2X1 XOR2_190 (.Y(N743),.A(N77),.B(N711));
XOR2X1 XOR2_191 (.Y(N744),.A(N81),.B(N712));
XOR2X1 XOR2_192 (.Y(N745),.A(N85),.B(N713));
XOR2X1 XOR2_193 (.Y(N746),.A(N89),.B(N714));
XOR2X1 XOR2_194 (.Y(N747),.A(N93),.B(N715));
XOR2X1 XOR2_195 (.Y(N748),.A(N97),.B(N716));
XOR2X1 XOR2_196 (.Y(N749),.A(N101),.B(N717));
XOR2X1 XOR2_197 (.Y(N750),.A(N105),.B(N718));
XOR2X1 XOR2_198 (.Y(N751),.A(N109),.B(N719));
XOR2X1 XOR2_199 (.Y(N752),.A(N113),.B(N720));
XOR2X1 XOR2_200 (.Y(N753),.A(N117),.B(N721));
XOR2X1 XOR2_201 (.Y(N754),.A(N121),.B(N722));
XOR2X1 XOR2_202 (.Y(N755),.A(N125),.B(N723));
endmodule