module c880 (N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,N219,N228,N237,N246,N255,N259,N260,N261,N267,N268,N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,N865,N866,N874,N878,N879,N880);
input N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,N219,N228,N237,N246,N255,N259,N260,N261,N267,N268;
output N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,N865,N866,N874,N878,N879,N880;
wire N269,N270,N273,N276,N279,N280,N284,N285,N286,N287,N290,N291,N292,N293,N294,N295,N296,N297,N298,N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N316,N317,N318,N319,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,N360,N363,N366,N369,N375,N376,N379,N382,N385,N392,N393,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N424,N425,N426,N427,N432,N437,N442,N443,N444,N445,N451,N460,N463,N466,N475,N476,N477,N478,N479,N480,N481,N482,N483,N488,N489,N490,N491,N492,N495,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N533,N536,N537,N538,N539,N540,N541,N542,N543,N544,N547,N550,N551,N552,N553,N557,N561,N565,N569,N573,N577,N581,N585,N586,N587,N588,N589,N590,N593,N596,N597,N600,N605,N606,N609,N615,N616,N619,N624,N625,N628,N631,N632,N635,N640,N641,N644,N650,N651,N654,N659,N660,N661,N662,N665,N669,N670,N673,N677,N678,N682,N686,N687,N692,N696,N697,N700,N704,N705,N708,N712,N713,N717,N721,N722,N727,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,N769,N770,N771,N772,N773,N777,N778,N781,N782,N785,N786,N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,N802,N803,N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N819,N822,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N851,N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,N867,N868,N869,N870,N871,N872,N873,N875,N876,N877;
AND2X1 AND_tmp1 (.Y(ttmp1),.A(N13),.B(N17));
AND2X1 AND_tmp2 (.Y(ttmp2),.A(N1),.B(ttmp1));
NAND2X1 NAND_tmp3 (.Y(N269),.A(N8),.B(ttmp2));
AND2X1 AND_tmp4 (.Y(ttmp4),.A(N13),.B(N17));
AND2X1 AND_tmp5 (.Y(ttmp5),.A(N1),.B(ttmp4));
NAND2X1 NAND_tmp6 (.Y(N270),.A(N26),.B(ttmp5));
AND2X1 AND_tmp7 (.Y(ttmp7),.A(N36),.B(N42));
AND2X1 AND_tmp8 (.Y(N273),.A(N29),.B(ttmp7));
AND2X1 AND_tmp9 (.Y(ttmp9),.A(N26),.B(N51));
AND2X1 AND_tmp10 (.Y(N276),.A(N1),.B(ttmp9));
AND2X1 AND_tmp11 (.Y(ttmp11),.A(N51),.B(N17));
AND2X1 AND_tmp12 (.Y(ttmp12),.A(N1),.B(ttmp11));
NAND2X1 NAND_tmp13 (.Y(N279),.A(N8),.B(ttmp12));
AND2X1 AND_tmp14 (.Y(ttmp14),.A(N13),.B(N55));
AND2X1 AND_tmp15 (.Y(ttmp15),.A(N1),.B(ttmp14));
NAND2X1 NAND_tmp16 (.Y(N280),.A(N8),.B(ttmp15));
AND2X1 AND_tmp17 (.Y(ttmp17),.A(N68),.B(N72));
AND2X1 AND_tmp18 (.Y(ttmp18),.A(N59),.B(ttmp17));
NAND2X1 NAND_tmp19 (.Y(N284),.A(N42),.B(ttmp18));
NAND2X1 NAND2_8 (.Y(N285),.A(N29),.B(N68));
AND2X1 AND_tmp20 (.Y(ttmp20),.A(N68),.B(N74));
NAND2X1 NAND_tmp21 (.Y(N286),.A(N59),.B(ttmp20));
AND2X1 AND_tmp22 (.Y(ttmp22),.A(N75),.B(N80));
AND2X1 AND_tmp23 (.Y(N287),.A(N29),.B(ttmp22));
AND2X1 AND_tmp24 (.Y(ttmp24),.A(N75),.B(N42));
AND2X1 AND_tmp25 (.Y(N290),.A(N29),.B(ttmp24));
AND2X1 AND_tmp26 (.Y(ttmp26),.A(N36),.B(N80));
AND2X1 AND_tmp27 (.Y(N291),.A(N29),.B(ttmp26));
AND2X1 AND_tmp28 (.Y(ttmp28),.A(N36),.B(N42));
AND2X1 AND_tmp29 (.Y(N292),.A(N29),.B(ttmp28));
AND2X1 AND_tmp30 (.Y(ttmp30),.A(N75),.B(N80));
AND2X1 AND_tmp31 (.Y(N293),.A(N59),.B(ttmp30));
AND2X1 AND_tmp32 (.Y(ttmp32),.A(N75),.B(N42));
AND2X1 AND_tmp33 (.Y(N294),.A(N59),.B(ttmp32));
AND2X1 AND_tmp34 (.Y(ttmp34),.A(N36),.B(N80));
AND2X1 AND_tmp35 (.Y(N295),.A(N59),.B(ttmp34));
AND2X1 AND_tmp36 (.Y(ttmp36),.A(N36),.B(N42));
AND2X1 AND_tmp37 (.Y(N296),.A(N59),.B(ttmp36));
AND2X1 AND2_18 (.Y(N297),.A(N85),.B(N86));
OR2X1 OR2_19 (.Y(N298),.A(N87),.B(N88));
NAND2X1 NAND2_20 (.Y(N301),.A(N91),.B(N96));
OR2X1 OR2_21 (.Y(N302),.A(N91),.B(N96));
NAND2X1 NAND2_22 (.Y(N303),.A(N101),.B(N106));
OR2X1 OR2_23 (.Y(N304),.A(N101),.B(N106));
NAND2X1 NAND2_24 (.Y(N305),.A(N111),.B(N116));
OR2X1 OR2_25 (.Y(N306),.A(N111),.B(N116));
NAND2X1 NAND2_26 (.Y(N307),.A(N121),.B(N126));
OR2X1 OR2_27 (.Y(N308),.A(N121),.B(N126));
AND2X1 AND2_28 (.Y(N309),.A(N8),.B(N138));
INVX1 NOT1_29 (.Y(N310),.A(N268));
AND2X1 AND2_30 (.Y(N316),.A(N51),.B(N138));
AND2X1 AND2_31 (.Y(N317),.A(N17),.B(N138));
AND2X1 AND2_32 (.Y(N318),.A(N152),.B(N138));
NAND2X1 NAND2_33 (.Y(N319),.A(N59),.B(N156));
NOR2X1 NOR2_34 (.Y(N322),.A(N17),.B(N42));
AND2X1 AND2_35 (.Y(N323),.A(N17),.B(N42));
NAND2X1 NAND2_36 (.Y(N324),.A(N159),.B(N165));
OR2X1 OR2_37 (.Y(N325),.A(N159),.B(N165));
NAND2X1 NAND2_38 (.Y(N326),.A(N171),.B(N177));
OR2X1 OR2_39 (.Y(N327),.A(N171),.B(N177));
NAND2X1 NAND2_40 (.Y(N328),.A(N183),.B(N189));
OR2X1 OR2_41 (.Y(N329),.A(N183),.B(N189));
NAND2X1 NAND2_42 (.Y(N330),.A(N195),.B(N201));
OR2X1 OR2_43 (.Y(N331),.A(N195),.B(N201));
AND2X1 AND2_44 (.Y(N332),.A(N210),.B(N91));
AND2X1 AND2_45 (.Y(N333),.A(N210),.B(N96));
AND2X1 AND2_46 (.Y(N334),.A(N210),.B(N101));
AND2X1 AND2_47 (.Y(N335),.A(N210),.B(N106));
AND2X1 AND2_48 (.Y(N336),.A(N210),.B(N111));
AND2X1 AND2_49 (.Y(N337),.A(N255),.B(N259));
AND2X1 AND2_50 (.Y(N338),.A(N210),.B(N116));
AND2X1 AND2_51 (.Y(N339),.A(N255),.B(N260));
AND2X1 AND2_52 (.Y(N340),.A(N210),.B(N121));
AND2X1 AND2_53 (.Y(N341),.A(N255),.B(N267));
INVX1 NOT1_54 (.Y(N342),.A(N269));
INVX1 NOT1_55 (.Y(N343),.A(N273));
OR2X1 OR2_56 (.Y(N344),.A(N270),.B(N273));
INVX1 NOT1_57 (.Y(N345),.A(N276));
INVX1 NOT1_58 (.Y(N346),.A(N276));
INVX1 NOT1_59 (.Y(N347),.A(N279));
NOR2X1 NOR2_60 (.Y(N348),.A(N280),.B(N284));
OR2X1 OR2_61 (.Y(N349),.A(N280),.B(N285));
OR2X1 OR2_62 (.Y(N350),.A(N280),.B(N286));
INVX1 NOT1_63 (.Y(N351),.A(N293));
INVX1 NOT1_64 (.Y(N352),.A(N294));
INVX1 NOT1_65 (.Y(N353),.A(N295));
INVX1 NOT1_66 (.Y(N354),.A(N296));
NAND2X1 NAND2_67 (.Y(N355),.A(N89),.B(N298));
AND2X1 AND2_68 (.Y(N356),.A(N90),.B(N298));
NAND2X1 NAND2_69 (.Y(N357),.A(N301),.B(N302));
NAND2X1 NAND2_70 (.Y(N360),.A(N303),.B(N304));
NAND2X1 NAND2_71 (.Y(N363),.A(N305),.B(N306));
NAND2X1 NAND2_72 (.Y(N366),.A(N307),.B(N308));
INVX1 NOT1_73 (.Y(N369),.A(N310));
NOR2X1 NOR2_74 (.Y(N375),.A(N322),.B(N323));
NAND2X1 NAND2_75 (.Y(N376),.A(N324),.B(N325));
NAND2X1 NAND2_76 (.Y(N379),.A(N326),.B(N327));
NAND2X1 NAND2_77 (.Y(N382),.A(N328),.B(N329));
NAND2X1 NAND2_78 (.Y(N385),.A(N330),.B(N331));
BUFX1 BUFF1_79 (.Y(N388),.A(N290));
BUFX1 BUFF1_80 (.Y(N389),.A(N291));
BUFX1 BUFF1_81 (.Y(N390),.A(N292));
BUFX1 BUFF1_82 (.Y(N391),.A(N297));
OR2X1 OR2_83 (.Y(N392),.A(N270),.B(N343));
INVX1 NOT1_84 (.Y(N393),.A(N345));
INVX1 NOT1_85 (.Y(N399),.A(N346));
AND2X1 AND2_86 (.Y(N400),.A(N348),.B(N73));
INVX1 NOT1_87 (.Y(N401),.A(N349));
INVX1 NOT1_88 (.Y(N402),.A(N350));
INVX1 NOT1_89 (.Y(N403),.A(N355));
INVX1 NOT1_90 (.Y(N404),.A(N357));
INVX1 NOT1_91 (.Y(N405),.A(N360));
AND2X1 AND2_92 (.Y(N406),.A(N357),.B(N360));
INVX1 NOT1_93 (.Y(N407),.A(N363));
INVX1 NOT1_94 (.Y(N408),.A(N366));
AND2X1 AND2_95 (.Y(N409),.A(N363),.B(N366));
NAND2X1 NAND2_96 (.Y(N410),.A(N347),.B(N352));
INVX1 NOT1_97 (.Y(N411),.A(N376));
INVX1 NOT1_98 (.Y(N412),.A(N379));
AND2X1 AND2_99 (.Y(N413),.A(N376),.B(N379));
INVX1 NOT1_100 (.Y(N414),.A(N382));
INVX1 NOT1_101 (.Y(N415),.A(N385));
AND2X1 AND2_102 (.Y(N416),.A(N382),.B(N385));
AND2X1 AND2_103 (.Y(N417),.A(N210),.B(N369));
BUFX1 BUFF1_104 (.Y(N418),.A(N342));
BUFX1 BUFF1_105 (.Y(N419),.A(N344));
BUFX1 BUFF1_106 (.Y(N420),.A(N351));
BUFX1 BUFF1_107 (.Y(N421),.A(N353));
BUFX1 BUFF1_108 (.Y(N422),.A(N354));
BUFX1 BUFF1_109 (.Y(N423),.A(N356));
INVX1 NOT1_110 (.Y(N424),.A(N400));
AND2X1 AND2_111 (.Y(N425),.A(N404),.B(N405));
AND2X1 AND2_112 (.Y(N426),.A(N407),.B(N408));
AND2X1 AND_tmp38 (.Y(ttmp38),.A(N393),.B(N55));
AND2X1 AND_tmp39 (.Y(N427),.A(N319),.B(ttmp38));
AND2X1 AND_tmp40 (.Y(ttmp40),.A(N17),.B(N287));
AND2X1 AND_tmp41 (.Y(N432),.A(N393),.B(ttmp40));
AND2X1 AND_tmp42 (.Y(ttmp42),.A(N287),.B(N55));
NAND2X1 NAND_tmp43 (.Y(N437),.A(N393),.B(ttmp42));
AND2X1 AND_tmp44 (.Y(ttmp44),.A(N156),.B(N393));
AND2X1 AND_tmp45 (.Y(ttmp45),.A(N375),.B(ttmp44));
NAND2X1 NAND_tmp46 (.Y(N442),.A(N59),.B(ttmp45));
AND2X1 AND_tmp47 (.Y(ttmp47),.A(N319),.B(N17));
NAND2X1 NAND_tmp48 (.Y(N443),.A(N393),.B(ttmp47));
AND2X1 AND2_118 (.Y(N444),.A(N411),.B(N412));
AND2X1 AND2_119 (.Y(N445),.A(N414),.B(N415));
BUFX1 BUFF1_120 (.Y(N446),.A(N392));
BUFX1 BUFF1_121 (.Y(N447),.A(N399));
BUFX1 BUFF1_122 (.Y(N448),.A(N401));
BUFX1 BUFF1_123 (.Y(N449),.A(N402));
BUFX1 BUFF1_124 (.Y(N450),.A(N403));
INVX1 NOT1_125 (.Y(N451),.A(N424));
NOR2X1 NOR2_126 (.Y(N460),.A(N406),.B(N425));
NOR2X1 NOR2_127 (.Y(N463),.A(N409),.B(N426));
NAND2X1 NAND2_128 (.Y(N466),.A(N442),.B(N410));
AND2X1 AND2_129 (.Y(N475),.A(N143),.B(N427));
AND2X1 AND2_130 (.Y(N476),.A(N310),.B(N432));
AND2X1 AND2_131 (.Y(N477),.A(N146),.B(N427));
AND2X1 AND2_132 (.Y(N478),.A(N310),.B(N432));
AND2X1 AND2_133 (.Y(N479),.A(N149),.B(N427));
AND2X1 AND2_134 (.Y(N480),.A(N310),.B(N432));
AND2X1 AND2_135 (.Y(N481),.A(N153),.B(N427));
AND2X1 AND2_136 (.Y(N482),.A(N310),.B(N432));
NAND2X1 NAND2_137 (.Y(N483),.A(N443),.B(N1));
OR2X1 OR2_138 (.Y(N488),.A(N369),.B(N437));
OR2X1 OR2_139 (.Y(N489),.A(N369),.B(N437));
OR2X1 OR2_140 (.Y(N490),.A(N369),.B(N437));
OR2X1 OR2_141 (.Y(N491),.A(N369),.B(N437));
NOR2X1 NOR2_142 (.Y(N492),.A(N413),.B(N444));
NOR2X1 NOR2_143 (.Y(N495),.A(N416),.B(N445));
NAND2X1 NAND2_144 (.Y(N498),.A(N130),.B(N460));
OR2X1 OR2_145 (.Y(N499),.A(N130),.B(N460));
NAND2X1 NAND2_146 (.Y(N500),.A(N463),.B(N135));
OR2X1 OR2_147 (.Y(N501),.A(N463),.B(N135));
AND2X1 AND2_148 (.Y(N502),.A(N91),.B(N466));
NOR2X1 NOR2_149 (.Y(N503),.A(N475),.B(N476));
AND2X1 AND2_150 (.Y(N504),.A(N96),.B(N466));
NOR2X1 NOR2_151 (.Y(N505),.A(N477),.B(N478));
AND2X1 AND2_152 (.Y(N506),.A(N101),.B(N466));
NOR2X1 NOR2_153 (.Y(N507),.A(N479),.B(N480));
AND2X1 AND2_154 (.Y(N508),.A(N106),.B(N466));
NOR2X1 NOR2_155 (.Y(N509),.A(N481),.B(N482));
AND2X1 AND2_156 (.Y(N510),.A(N143),.B(N483));
AND2X1 AND2_157 (.Y(N511),.A(N111),.B(N466));
AND2X1 AND2_158 (.Y(N512),.A(N146),.B(N483));
AND2X1 AND2_159 (.Y(N513),.A(N116),.B(N466));
AND2X1 AND2_160 (.Y(N514),.A(N149),.B(N483));
AND2X1 AND2_161 (.Y(N515),.A(N121),.B(N466));
AND2X1 AND2_162 (.Y(N516),.A(N153),.B(N483));
AND2X1 AND2_163 (.Y(N517),.A(N126),.B(N466));
NAND2X1 NAND2_164 (.Y(N518),.A(N130),.B(N492));
OR2X1 OR2_165 (.Y(N519),.A(N130),.B(N492));
NAND2X1 NAND2_166 (.Y(N520),.A(N495),.B(N207));
OR2X1 OR2_167 (.Y(N521),.A(N495),.B(N207));
AND2X1 AND2_168 (.Y(N522),.A(N451),.B(N159));
AND2X1 AND2_169 (.Y(N523),.A(N451),.B(N165));
AND2X1 AND2_170 (.Y(N524),.A(N451),.B(N171));
AND2X1 AND2_171 (.Y(N525),.A(N451),.B(N177));
AND2X1 AND2_172 (.Y(N526),.A(N451),.B(N183));
NAND2X1 NAND2_173 (.Y(N527),.A(N451),.B(N189));
NAND2X1 NAND2_174 (.Y(N528),.A(N451),.B(N195));
NAND2X1 NAND2_175 (.Y(N529),.A(N451),.B(N201));
NAND2X1 NAND2_176 (.Y(N530),.A(N498),.B(N499));
NAND2X1 NAND2_177 (.Y(N533),.A(N500),.B(N501));
NOR2X1 NOR2_178 (.Y(N536),.A(N309),.B(N502));
NOR2X1 NOR2_179 (.Y(N537),.A(N316),.B(N504));
NOR2X1 NOR2_180 (.Y(N538),.A(N317),.B(N506));
NOR2X1 NOR2_181 (.Y(N539),.A(N318),.B(N508));
NOR2X1 NOR2_182 (.Y(N540),.A(N510),.B(N511));
NOR2X1 NOR2_183 (.Y(N541),.A(N512),.B(N513));
NOR2X1 NOR2_184 (.Y(N542),.A(N514),.B(N515));
NOR2X1 NOR2_185 (.Y(N543),.A(N516),.B(N517));
NAND2X1 NAND2_186 (.Y(N544),.A(N518),.B(N519));
NAND2X1 NAND2_187 (.Y(N547),.A(N520),.B(N521));
INVX1 NOT1_188 (.Y(N550),.A(N530));
INVX1 NOT1_189 (.Y(N551),.A(N533));
AND2X1 AND2_190 (.Y(N552),.A(N530),.B(N533));
NAND2X1 NAND2_191 (.Y(N553),.A(N536),.B(N503));
NAND2X1 NAND2_192 (.Y(N557),.A(N537),.B(N505));
NAND2X1 NAND2_193 (.Y(N561),.A(N538),.B(N507));
NAND2X1 NAND2_194 (.Y(N565),.A(N539),.B(N509));
NAND2X1 NAND2_195 (.Y(N569),.A(N488),.B(N540));
NAND2X1 NAND2_196 (.Y(N573),.A(N489),.B(N541));
NAND2X1 NAND2_197 (.Y(N577),.A(N490),.B(N542));
NAND2X1 NAND2_198 (.Y(N581),.A(N491),.B(N543));
INVX1 NOT1_199 (.Y(N585),.A(N544));
INVX1 NOT1_200 (.Y(N586),.A(N547));
AND2X1 AND2_201 (.Y(N587),.A(N544),.B(N547));
AND2X1 AND2_202 (.Y(N588),.A(N550),.B(N551));
AND2X1 AND2_203 (.Y(N589),.A(N585),.B(N586));
NAND2X1 NAND2_204 (.Y(N590),.A(N553),.B(N159));
OR2X1 OR2_205 (.Y(N593),.A(N553),.B(N159));
AND2X1 AND2_206 (.Y(N596),.A(N246),.B(N553));
NAND2X1 NAND2_207 (.Y(N597),.A(N557),.B(N165));
OR2X1 OR2_208 (.Y(N600),.A(N557),.B(N165));
AND2X1 AND2_209 (.Y(N605),.A(N246),.B(N557));
NAND2X1 NAND2_210 (.Y(N606),.A(N561),.B(N171));
OR2X1 OR2_211 (.Y(N609),.A(N561),.B(N171));
AND2X1 AND2_212 (.Y(N615),.A(N246),.B(N561));
NAND2X1 NAND2_213 (.Y(N616),.A(N565),.B(N177));
OR2X1 OR2_214 (.Y(N619),.A(N565),.B(N177));
AND2X1 AND2_215 (.Y(N624),.A(N246),.B(N565));
NAND2X1 NAND2_216 (.Y(N625),.A(N569),.B(N183));
OR2X1 OR2_217 (.Y(N628),.A(N569),.B(N183));
AND2X1 AND2_218 (.Y(N631),.A(N246),.B(N569));
NAND2X1 NAND2_219 (.Y(N632),.A(N573),.B(N189));
OR2X1 OR2_220 (.Y(N635),.A(N573),.B(N189));
AND2X1 AND2_221 (.Y(N640),.A(N246),.B(N573));
NAND2X1 NAND2_222 (.Y(N641),.A(N577),.B(N195));
OR2X1 OR2_223 (.Y(N644),.A(N577),.B(N195));
AND2X1 AND2_224 (.Y(N650),.A(N246),.B(N577));
NAND2X1 NAND2_225 (.Y(N651),.A(N581),.B(N201));
OR2X1 OR2_226 (.Y(N654),.A(N581),.B(N201));
AND2X1 AND2_227 (.Y(N659),.A(N246),.B(N581));
NOR2X1 NOR2_228 (.Y(N660),.A(N552),.B(N588));
NOR2X1 NOR2_229 (.Y(N661),.A(N587),.B(N589));
INVX1 NOT1_230 (.Y(N662),.A(N590));
AND2X1 AND2_231 (.Y(N665),.A(N593),.B(N590));
NOR2X1 NOR2_232 (.Y(N669),.A(N596),.B(N522));
INVX1 NOT1_233 (.Y(N670),.A(N597));
AND2X1 AND2_234 (.Y(N673),.A(N600),.B(N597));
NOR2X1 NOR2_235 (.Y(N677),.A(N605),.B(N523));
INVX1 NOT1_236 (.Y(N678),.A(N606));
AND2X1 AND2_237 (.Y(N682),.A(N609),.B(N606));
NOR2X1 NOR2_238 (.Y(N686),.A(N615),.B(N524));
INVX1 NOT1_239 (.Y(N687),.A(N616));
AND2X1 AND2_240 (.Y(N692),.A(N619),.B(N616));
NOR2X1 NOR2_241 (.Y(N696),.A(N624),.B(N525));
INVX1 NOT1_242 (.Y(N697),.A(N625));
AND2X1 AND2_243 (.Y(N700),.A(N628),.B(N625));
NOR2X1 NOR2_244 (.Y(N704),.A(N631),.B(N526));
INVX1 NOT1_245 (.Y(N705),.A(N632));
AND2X1 AND2_246 (.Y(N708),.A(N635),.B(N632));
NOR2X1 NOR2_247 (.Y(N712),.A(N337),.B(N640));
INVX1 NOT1_248 (.Y(N713),.A(N641));
AND2X1 AND2_249 (.Y(N717),.A(N644),.B(N641));
NOR2X1 NOR2_250 (.Y(N721),.A(N339),.B(N650));
INVX1 NOT1_251 (.Y(N722),.A(N651));
AND2X1 AND2_252 (.Y(N727),.A(N654),.B(N651));
NOR2X1 NOR2_253 (.Y(N731),.A(N341),.B(N659));
NAND2X1 NAND2_254 (.Y(N732),.A(N654),.B(N261));
AND2X1 AND_tmp49 (.Y(ttmp49),.A(N654),.B(N261));
NAND2X1 NAND_tmp50 (.Y(N733),.A(N644),.B(ttmp49));
AND2X1 AND_tmp51 (.Y(ttmp51),.A(N654),.B(N261));
AND2X1 AND_tmp52 (.Y(ttmp52),.A(N635),.B(ttmp51));
NAND2X1 NAND_tmp53 (.Y(N734),.A(N644),.B(ttmp52));
INVX1 NOT1_257 (.Y(N735),.A(N662));
AND2X1 AND2_258 (.Y(N736),.A(N228),.B(N665));
AND2X1 AND2_259 (.Y(N737),.A(N237),.B(N662));
INVX1 NOT1_260 (.Y(N738),.A(N670));
AND2X1 AND2_261 (.Y(N739),.A(N228),.B(N673));
AND2X1 AND2_262 (.Y(N740),.A(N237),.B(N670));
INVX1 NOT1_263 (.Y(N741),.A(N678));
AND2X1 AND2_264 (.Y(N742),.A(N228),.B(N682));
AND2X1 AND2_265 (.Y(N743),.A(N237),.B(N678));
INVX1 NOT1_266 (.Y(N744),.A(N687));
AND2X1 AND2_267 (.Y(N745),.A(N228),.B(N692));
AND2X1 AND2_268 (.Y(N746),.A(N237),.B(N687));
INVX1 NOT1_269 (.Y(N747),.A(N697));
AND2X1 AND2_270 (.Y(N748),.A(N228),.B(N700));
AND2X1 AND2_271 (.Y(N749),.A(N237),.B(N697));
INVX1 NOT1_272 (.Y(N750),.A(N705));
AND2X1 AND2_273 (.Y(N751),.A(N228),.B(N708));
AND2X1 AND2_274 (.Y(N752),.A(N237),.B(N705));
INVX1 NOT1_275 (.Y(N753),.A(N713));
AND2X1 AND2_276 (.Y(N754),.A(N228),.B(N717));
AND2X1 AND2_277 (.Y(N755),.A(N237),.B(N713));
INVX1 NOT1_278 (.Y(N756),.A(N722));
NOR2X1 NOR2_279 (.Y(N757),.A(N727),.B(N261));
AND2X1 AND2_280 (.Y(N758),.A(N727),.B(N261));
AND2X1 AND2_281 (.Y(N759),.A(N228),.B(N727));
AND2X1 AND2_282 (.Y(N760),.A(N237),.B(N722));
NAND2X1 NAND2_283 (.Y(N761),.A(N644),.B(N722));
NAND2X1 NAND2_284 (.Y(N762),.A(N635),.B(N713));
AND2X1 AND_tmp54 (.Y(ttmp54),.A(N644),.B(N722));
NAND2X1 NAND_tmp55 (.Y(N763),.A(N635),.B(ttmp54));
NAND2X1 NAND2_286 (.Y(N764),.A(N609),.B(N687));
NAND2X1 NAND2_287 (.Y(N765),.A(N600),.B(N678));
AND2X1 AND_tmp56 (.Y(ttmp56),.A(N609),.B(N687));
NAND2X1 NAND_tmp57 (.Y(N766),.A(N600),.B(ttmp56));
BUFX1 BUFF1_289 (.Y(N767),.A(N660));
BUFX1 BUFF1_290 (.Y(N768),.A(N661));
NOR2X1 NOR2_291 (.Y(N769),.A(N736),.B(N737));
NOR2X1 NOR2_292 (.Y(N770),.A(N739),.B(N740));
NOR2X1 NOR2_293 (.Y(N771),.A(N742),.B(N743));
NOR2X1 NOR2_294 (.Y(N772),.A(N745),.B(N746));
AND2X1 AND_tmp58 (.Y(ttmp58),.A(N763),.B(N734));
AND2X1 AND_tmp59 (.Y(ttmp59),.A(N750),.B(ttmp58));
NAND2X1 NAND_tmp60 (.Y(N773),.A(N762),.B(ttmp59));
NOR2X1 NOR2_296 (.Y(N777),.A(N748),.B(N749));
AND2X1 AND_tmp61 (.Y(ttmp61),.A(N761),.B(N733));
NAND2X1 NAND_tmp62 (.Y(N778),.A(N753),.B(ttmp61));
NOR2X1 NOR2_298 (.Y(N781),.A(N751),.B(N752));
NAND2X1 NAND2_299 (.Y(N782),.A(N756),.B(N732));
NOR2X1 NOR2_300 (.Y(N785),.A(N754),.B(N755));
NOR2X1 NOR2_301 (.Y(N786),.A(N757),.B(N758));
NOR2X1 NOR2_302 (.Y(N787),.A(N759),.B(N760));
NOR2X1 NOR2_303 (.Y(N788),.A(N700),.B(N773));
AND2X1 AND2_304 (.Y(N789),.A(N700),.B(N773));
NOR2X1 NOR2_305 (.Y(N790),.A(N708),.B(N778));
AND2X1 AND2_306 (.Y(N791),.A(N708),.B(N778));
NOR2X1 NOR2_307 (.Y(N792),.A(N717),.B(N782));
AND2X1 AND2_308 (.Y(N793),.A(N717),.B(N782));
AND2X1 AND2_309 (.Y(N794),.A(N219),.B(N786));
NAND2X1 NAND2_310 (.Y(N795),.A(N628),.B(N773));
NAND2X1 NAND2_311 (.Y(N796),.A(N795),.B(N747));
NOR2X1 NOR2_312 (.Y(N802),.A(N788),.B(N789));
NOR2X1 NOR2_313 (.Y(N803),.A(N790),.B(N791));
NOR2X1 NOR2_314 (.Y(N804),.A(N792),.B(N793));
NOR2X1 NOR2_315 (.Y(N805),.A(N340),.B(N794));
NOR2X1 NOR2_316 (.Y(N806),.A(N692),.B(N796));
AND2X1 AND2_317 (.Y(N807),.A(N692),.B(N796));
AND2X1 AND2_318 (.Y(N808),.A(N219),.B(N802));
AND2X1 AND2_319 (.Y(N809),.A(N219),.B(N803));
AND2X1 AND2_320 (.Y(N810),.A(N219),.B(N804));
AND2X1 AND_tmp63 (.Y(ttmp63),.A(N731),.B(N529));
AND2X1 AND_tmp64 (.Y(ttmp64),.A(N805),.B(ttmp63));
NAND2X1 NAND_tmp65 (.Y(N811),.A(N787),.B(ttmp64));
NAND2X1 NAND2_322 (.Y(N812),.A(N619),.B(N796));
AND2X1 AND_tmp66 (.Y(ttmp66),.A(N619),.B(N796));
NAND2X1 NAND_tmp67 (.Y(N813),.A(N609),.B(ttmp66));
AND2X1 AND_tmp68 (.Y(ttmp68),.A(N619),.B(N796));
AND2X1 AND_tmp69 (.Y(ttmp69),.A(N600),.B(ttmp68));
NAND2X1 NAND_tmp70 (.Y(N814),.A(N609),.B(ttmp69));
AND2X1 AND_tmp71 (.Y(ttmp71),.A(N766),.B(N814));
AND2X1 AND_tmp72 (.Y(ttmp72),.A(N738),.B(ttmp71));
NAND2X1 NAND_tmp73 (.Y(N815),.A(N765),.B(ttmp72));
AND2X1 AND_tmp74 (.Y(ttmp74),.A(N764),.B(N813));
NAND2X1 NAND_tmp75 (.Y(N819),.A(N741),.B(ttmp74));
NAND2X1 NAND2_327 (.Y(N822),.A(N744),.B(N812));
NOR2X1 NOR2_328 (.Y(N825),.A(N806),.B(N807));
NOR2X1 NOR2_329 (.Y(N826),.A(N335),.B(N808));
NOR2X1 NOR2_330 (.Y(N827),.A(N336),.B(N809));
NOR2X1 NOR2_331 (.Y(N828),.A(N338),.B(N810));
INVX1 NOT1_332 (.Y(N829),.A(N811));
NOR2X1 NOR2_333 (.Y(N830),.A(N665),.B(N815));
AND2X1 AND2_334 (.Y(N831),.A(N665),.B(N815));
NOR2X1 NOR2_335 (.Y(N832),.A(N673),.B(N819));
AND2X1 AND2_336 (.Y(N833),.A(N673),.B(N819));
NOR2X1 NOR2_337 (.Y(N834),.A(N682),.B(N822));
AND2X1 AND2_338 (.Y(N835),.A(N682),.B(N822));
AND2X1 AND2_339 (.Y(N836),.A(N219),.B(N825));
AND2X1 AND_tmp76 (.Y(ttmp76),.A(N777),.B(N704));
NAND2X1 NAND_tmp77 (.Y(N837),.A(N826),.B(ttmp76));
AND2X1 AND_tmp78 (.Y(ttmp78),.A(N712),.B(N527));
AND2X1 AND_tmp79 (.Y(ttmp79),.A(N827),.B(ttmp78));
NAND2X1 NAND_tmp80 (.Y(N838),.A(N781),.B(ttmp79));
AND2X1 AND_tmp81 (.Y(ttmp81),.A(N721),.B(N528));
AND2X1 AND_tmp82 (.Y(ttmp82),.A(N828),.B(ttmp81));
NAND2X1 NAND_tmp83 (.Y(N839),.A(N785),.B(ttmp82));
INVX1 NOT1_343 (.Y(N840),.A(N829));
NAND2X1 NAND2_344 (.Y(N841),.A(N815),.B(N593));
NOR2X1 NOR2_345 (.Y(N842),.A(N830),.B(N831));
NOR2X1 NOR2_346 (.Y(N843),.A(N832),.B(N833));
NOR2X1 NOR2_347 (.Y(N844),.A(N834),.B(N835));
NOR2X1 NOR2_348 (.Y(N845),.A(N334),.B(N836));
INVX1 NOT1_349 (.Y(N846),.A(N837));
INVX1 NOT1_350 (.Y(N847),.A(N838));
INVX1 NOT1_351 (.Y(N848),.A(N839));
AND2X1 AND2_352 (.Y(N849),.A(N735),.B(N841));
BUFX1 BUFF1_353 (.Y(N850),.A(N840));
AND2X1 AND2_354 (.Y(N851),.A(N219),.B(N842));
AND2X1 AND2_355 (.Y(N852),.A(N219),.B(N843));
AND2X1 AND2_356 (.Y(N853),.A(N219),.B(N844));
AND2X1 AND_tmp84 (.Y(ttmp84),.A(N772),.B(N696));
NAND2X1 NAND_tmp85 (.Y(N854),.A(N845),.B(ttmp84));
INVX1 NOT1_358 (.Y(N855),.A(N846));
INVX1 NOT1_359 (.Y(N856),.A(N847));
INVX1 NOT1_360 (.Y(N857),.A(N848));
INVX1 NOT1_361 (.Y(N858),.A(N849));
NOR2X1 NOR2_362 (.Y(N859),.A(N417),.B(N851));
NOR2X1 NOR2_363 (.Y(N860),.A(N332),.B(N852));
NOR2X1 NOR2_364 (.Y(N861),.A(N333),.B(N853));
INVX1 NOT1_365 (.Y(N862),.A(N854));
BUFX1 BUFF1_366 (.Y(N863),.A(N855));
BUFX1 BUFF1_367 (.Y(N864),.A(N856));
BUFX1 BUFF1_368 (.Y(N865),.A(N857));
BUFX1 BUFF1_369 (.Y(N866),.A(N858));
AND2X1 AND_tmp86 (.Y(ttmp86),.A(N769),.B(N669));
NAND2X1 NAND_tmp87 (.Y(N867),.A(N859),.B(ttmp86));
AND2X1 AND_tmp88 (.Y(ttmp88),.A(N770),.B(N677));
NAND2X1 NAND_tmp89 (.Y(N868),.A(N860),.B(ttmp88));
AND2X1 AND_tmp90 (.Y(ttmp90),.A(N771),.B(N686));
NAND2X1 NAND_tmp91 (.Y(N869),.A(N861),.B(ttmp90));
INVX1 NOT1_373 (.Y(N870),.A(N862));
INVX1 NOT1_374 (.Y(N871),.A(N867));
INVX1 NOT1_375 (.Y(N872),.A(N868));
INVX1 NOT1_376 (.Y(N873),.A(N869));
BUFX1 BUFF1_377 (.Y(N874),.A(N870));
INVX1 NOT1_378 (.Y(N875),.A(N871));
INVX1 NOT1_379 (.Y(N876),.A(N872));
INVX1 NOT1_380 (.Y(N877),.A(N873));
BUFX1 BUFF1_381 (.Y(N878),.A(N875));
BUFX1 BUFF1_382 (.Y(N879),.A(N876));
BUFX1 BUFF1_383 (.Y(N880),.A(N877));
endmodule