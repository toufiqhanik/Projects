.Option ingold=2 accurate
.OPTION MEASDGT=8
.OPTION NUMDGT=10
+ RUNLVL=5 ACCURATE
.op
.PARAM LMIN='50E-9'
.PARAM VDD_VALUE=1.2
.PARAM VDD_HALF=0.6
.OPTION BRIEF=1

.OPTION POST=2
.OPTION MEASFORM=3
.OPTION PROBE=1
***fast
.option NOTOP NOELCHK
.option AUTOSTOP
*****
VSUPPLY VDD1 0 VDD_VALUE
Rres1 VDD1 VDD 50
VSUPPLYGND GND 0 0

.include './trans_model_nk'
.include './all_gates_anik'
.temp 25

.TRAN 10p 142N START=0N

*Vinputclk CLK PULSE (V1 V2 Td Tr Tf Pw Period)
Vinputclk CLK GND PULSE (0V 1.2V 5ns 0.001ns 0.001ns 5ns 10ns)
Vinputrstn RSTn GND PWL(0 0 9.999n 0 10n VDD_VALUE)
VinputDrdy Drdy GND PWL(0 0 19.999n 0 20n VDD_VALUE)
VinputKrdy Krdy GND PWL(0 0 9.999n 0 10n VDD_VALUE 19.999n VDD_VALUE 20n 0)

VinputEnDec EncDec GND PWL(0 0)
VinputEn EN GND PWL(0 VDD_VALUE)


paramvar


xAES_Comp_ENCa/BSYrg_reg n8244 CLK BSY_E n981 VDD GND DFF_X1
xAES_Comp_ENCa/Rrg_reg_0 n8112 CLK \AES_Comp_ENCa/Rrg_0 n813 VDD GND DFF_X1
xAES_Comp_ENCa/Rrg_reg_1 n8109 CLK \AES_Comp_ENCa/Rrg_1 dummy1 VDD GND DFF_X1
xAES_Comp_ENCa/Rrg_reg_2 n8113 CLK \AES_Comp_ENCa/Rrg_2 dummy2 VDD GND DFF_X1
xAES_Comp_ENCa/Rrg_reg_3 n8108 CLK \AES_Comp_ENCa/Rrg_3 n814 VDD GND DFF_X1
xAES_Comp_ENCa/Rrg_reg_4 n8107 CLK \AES_Comp_ENCa/Rrg_4 n815 VDD GND DFF_X1
xAES_Comp_ENCa/Rrg_reg_5 n8106 CLK \AES_Comp_ENCa/Rrg_5 dummy3 VDD GND DFF_X1
xAES_Comp_ENCa/Rrg_reg_6 n8105 CLK \AES_Comp_ENCa/Rrg_6 dummy4 VDD GND DFF_X1
xAES_Comp_ENCa/Rrg_reg_7 n8104 CLK \AES_Comp_ENCa/Rrg_7 n816 VDD GND DFF_X1
xAES_Comp_ENCa/Rrg_reg_8 n8103 CLK \AES_Comp_ENCa/Rrg_8 dummy5 VDD GND DFF_X1
xAES_Comp_ENCa/Rrg_reg_9 n8102 CLK \AES_Comp_ENCa/Rrg_9 n817 VDD GND DFF_X1
xAES_Comp_ENCa/Kvldrg_reg n8242 CLK Kvld_E n818 VDD GND DFF_X1
xKvld_reg_reg n8241 CLK Kvld_reg dummy6 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_2 n8114 CLK \AES_Comp_ENCa/Krg_2 n683 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_3 n8115 CLK \AES_Comp_ENCa/Krg_3 n684 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_4 n8116 CLK \AES_Comp_ENCa/Krg_4 n685 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_5 n8117 CLK \AES_Comp_ENCa/Krg_5 n686 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_6 n8118 CLK \AES_Comp_ENCa/Krg_6 n687 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_7 n8119 CLK \AES_Comp_ENCa/Krg_7 n688 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_8 n8120 CLK \AES_Comp_ENCa/Krg_8 n689 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_9 n8121 CLK \AES_Comp_ENCa/Krg_9 n690 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_10 n8122 CLK \AES_Comp_ENCa/Krg_10 n691 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_11 n8123 CLK \AES_Comp_ENCa/Krg_11 n692 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_12 n8124 CLK \AES_Comp_ENCa/Krg_12 n693 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_13 n8125 CLK \AES_Comp_ENCa/Krg_13 n694 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_14 n8126 CLK \AES_Comp_ENCa/Krg_14 n695 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_15 n8127 CLK \AES_Comp_ENCa/Krg_15 n696 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_16 n8128 CLK \AES_Comp_ENCa/Krg_16 n697 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_17 n8129 CLK \AES_Comp_ENCa/Krg_17 n698 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_18 n8130 CLK \AES_Comp_ENCa/Krg_18 n699 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_19 n8131 CLK \AES_Comp_ENCa/Krg_19 n700 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_20 n8132 CLK \AES_Comp_ENCa/Krg_20 n701 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_21 n8133 CLK \AES_Comp_ENCa/Krg_21 n702 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_22 n8134 CLK \AES_Comp_ENCa/Krg_22 n703 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_23 n8135 CLK \AES_Comp_ENCa/Krg_23 n704 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_24 n8136 CLK \AES_Comp_ENCa/Krg_24 n705 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_25 n8137 CLK \AES_Comp_ENCa/Krg_25 n706 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_26 n8138 CLK \AES_Comp_ENCa/Krg_26 n707 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_27 n8139 CLK \AES_Comp_ENCa/Krg_27 n708 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_28 n8140 CLK \AES_Comp_ENCa/Krg_28 n709 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_29 n8141 CLK \AES_Comp_ENCa/Krg_29 n710 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_1 n8142 CLK \AES_Comp_ENCa/Krg_1 n682 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_30 n8143 CLK \AES_Comp_ENCa/Krg_30 n711 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_31 n8144 CLK \AES_Comp_ENCa/Krg_31 n712 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_32 n8145 CLK \AES_Comp_ENCa/Krg_32 n713 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_33 n8146 CLK \AES_Comp_ENCa/Krg_33 n714 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_34 n8147 CLK \AES_Comp_ENCa/Krg_34 n715 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_35 n8148 CLK \AES_Comp_ENCa/Krg_35 n716 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_36 n8149 CLK \AES_Comp_ENCa/Krg_36 n717 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_37 n8150 CLK \AES_Comp_ENCa/Krg_37 n718 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_38 n8151 CLK \AES_Comp_ENCa/Krg_38 n719 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_39 n8152 CLK \AES_Comp_ENCa/Krg_39 n720 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_40 n8153 CLK \AES_Comp_ENCa/Krg_40 n721 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_41 n8154 CLK \AES_Comp_ENCa/Krg_41 n722 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_42 n8155 CLK \AES_Comp_ENCa/Krg_42 n723 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_43 n8156 CLK \AES_Comp_ENCa/Krg_43 n724 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_44 n8157 CLK \AES_Comp_ENCa/Krg_44 n725 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_45 n8158 CLK \AES_Comp_ENCa/Krg_45 n726 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_46 n8159 CLK \AES_Comp_ENCa/Krg_46 n727 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_47 n8160 CLK \AES_Comp_ENCa/Krg_47 n728 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_48 n8161 CLK \AES_Comp_ENCa/Krg_48 n729 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_49 n8162 CLK \AES_Comp_ENCa/Krg_49 n730 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_50 n8163 CLK \AES_Comp_ENCa/Krg_50 n731 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_51 n8164 CLK \AES_Comp_ENCa/Krg_51 n732 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_52 n8165 CLK \AES_Comp_ENCa/Krg_52 n733 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_53 n8166 CLK \AES_Comp_ENCa/Krg_53 n734 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_54 n8167 CLK \AES_Comp_ENCa/Krg_54 n735 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_55 n8168 CLK \AES_Comp_ENCa/Krg_55 n736 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_56 n8169 CLK \AES_Comp_ENCa/Krg_56 n737 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_57 n8170 CLK \AES_Comp_ENCa/Krg_57 n738 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_58 n8171 CLK \AES_Comp_ENCa/Krg_58 n739 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_59 n8172 CLK \AES_Comp_ENCa/Krg_59 n740 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_60 n8173 CLK \AES_Comp_ENCa/Krg_60 n741 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_61 n8174 CLK \AES_Comp_ENCa/Krg_61 n742 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_62 n8175 CLK \AES_Comp_ENCa/Krg_62 n743 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_63 n8176 CLK \AES_Comp_ENCa/Krg_63 n744 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_64 n8177 CLK \AES_Comp_ENCa/Krg_64 n745 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_65 n8178 CLK \AES_Comp_ENCa/Krg_65 n746 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_66 n8179 CLK \AES_Comp_ENCa/Krg_66 n747 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_67 n8180 CLK \AES_Comp_ENCa/Krg_67 n748 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_68 n8181 CLK \AES_Comp_ENCa/Krg_68 n749 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_69 n8182 CLK \AES_Comp_ENCa/Krg_69 n750 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_70 n8183 CLK \AES_Comp_ENCa/Krg_70 n751 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_71 n8184 CLK \AES_Comp_ENCa/Krg_71 n752 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_72 n8185 CLK \AES_Comp_ENCa/Krg_72 n753 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_73 n8186 CLK \AES_Comp_ENCa/Krg_73 n754 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_74 n8187 CLK \AES_Comp_ENCa/Krg_74 n755 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_75 n8188 CLK \AES_Comp_ENCa/Krg_75 n756 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_76 n8189 CLK \AES_Comp_ENCa/Krg_76 n757 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_77 n8190 CLK \AES_Comp_ENCa/Krg_77 n758 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_78 n8191 CLK \AES_Comp_ENCa/Krg_78 n759 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_79 n8192 CLK \AES_Comp_ENCa/Krg_79 n760 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_80 n8193 CLK \AES_Comp_ENCa/Krg_80 n761 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_81 n8194 CLK \AES_Comp_ENCa/Krg_81 n762 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_82 n8195 CLK \AES_Comp_ENCa/Krg_82 n763 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_83 n8196 CLK \AES_Comp_ENCa/Krg_83 n764 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_84 n8197 CLK \AES_Comp_ENCa/Krg_84 n765 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_85 n8198 CLK \AES_Comp_ENCa/Krg_85 n766 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_86 n8199 CLK \AES_Comp_ENCa/Krg_86 n767 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_87 n8200 CLK \AES_Comp_ENCa/Krg_87 n768 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_88 n8201 CLK \AES_Comp_ENCa/Krg_88 n769 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_89 n8202 CLK \AES_Comp_ENCa/Krg_89 n770 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_90 n8203 CLK \AES_Comp_ENCa/Krg_90 n771 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_91 n8204 CLK \AES_Comp_ENCa/Krg_91 n772 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_92 n8205 CLK \AES_Comp_ENCa/Krg_92 n773 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_93 n8206 CLK \AES_Comp_ENCa/Krg_93 n774 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_94 n8207 CLK \AES_Comp_ENCa/Krg_94 n775 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_95 n8208 CLK \AES_Comp_ENCa/Krg_95 n776 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_96 n8209 CLK \AES_Comp_ENCa/Krg_96 n777 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_97 n8210 CLK \AES_Comp_ENCa/Krg_97 n778 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_98 n8211 CLK \AES_Comp_ENCa/Krg_98 n779 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_99 n8212 CLK \AES_Comp_ENCa/Krg_99 n780 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_100 n8213 CLK \AES_Comp_ENCa/Krg_100 n781 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_101 n8214 CLK \AES_Comp_ENCa/Krg_101 n782 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_102 n8215 CLK \AES_Comp_ENCa/Krg_102 n783 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_103 n8216 CLK \AES_Comp_ENCa/Krg_103 n784 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_104 n8217 CLK \AES_Comp_ENCa/Krg_104 n785 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_105 n8218 CLK \AES_Comp_ENCa/Krg_105 n786 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_106 n8219 CLK \AES_Comp_ENCa/Krg_106 n787 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_107 n8220 CLK \AES_Comp_ENCa/Krg_107 n788 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_108 n8221 CLK \AES_Comp_ENCa/Krg_108 n789 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_109 n8222 CLK \AES_Comp_ENCa/Krg_109 n790 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_110 n8223 CLK \AES_Comp_ENCa/Krg_110 n791 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_111 n8224 CLK \AES_Comp_ENCa/Krg_111 n792 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_112 n8225 CLK \AES_Comp_ENCa/Krg_112 n793 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_113 n8226 CLK \AES_Comp_ENCa/Krg_113 n794 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_114 n8227 CLK \AES_Comp_ENCa/Krg_114 n795 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_115 n8228 CLK \AES_Comp_ENCa/Krg_115 n796 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_116 n8229 CLK \AES_Comp_ENCa/Krg_116 n797 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_117 n8230 CLK \AES_Comp_ENCa/Krg_117 n798 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_118 n8231 CLK \AES_Comp_ENCa/Krg_118 n799 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_119 n8232 CLK \AES_Comp_ENCa/Krg_119 n800 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_120 n8233 CLK \AES_Comp_ENCa/Krg_120 n801 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_121 n8234 CLK \AES_Comp_ENCa/Krg_121 n802 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_122 n8235 CLK \AES_Comp_ENCa/Krg_122 n803 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_123 n8236 CLK \AES_Comp_ENCa/Krg_123 n804 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_124 n8237 CLK \AES_Comp_ENCa/Krg_124 n805 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_125 n8238 CLK \AES_Comp_ENCa/Krg_125 n806 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_126 n8239 CLK \AES_Comp_ENCa/Krg_126 n807 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_127 n8240 CLK \AES_Comp_ENCa/Krg_127 n808 VDD GND DFF_X1
xAES_Comp_ENCa/Krg_reg_0 n8243 CLK \AES_Comp_ENCa/Krg_0 n681 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_0 n8101 CLK \AES_Comp_ENCa/KrgX_0 n824 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_40 n8061 CLK \AES_Comp_ENCa/KrgX_40 n893 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_8 n8093 CLK \AES_Comp_ENCa/KrgX_8 n839 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_48 n8053 CLK \AES_Comp_ENCa/KrgX_48 n901 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_16 n8085 CLK \AES_Comp_ENCa/KrgX_16 n854 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_56 n8045 CLK \AES_Comp_ENCa/KrgX_56 n909 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_24 n8077 CLK \AES_Comp_ENCa/KrgX_24 n875 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_36 n8065 CLK \AES_Comp_ENCa/KrgX_36 n889 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_4 n8097 CLK \AES_Comp_ENCa/KrgX_4 n829 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_41 n8060 CLK \AES_Comp_ENCa/KrgX_41 n894 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_9 n8092 CLK \AES_Comp_ENCa/KrgX_9 n840 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_49 n8052 CLK \AES_Comp_ENCa/KrgX_49 n902 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_17 n8084 CLK \AES_Comp_ENCa/KrgX_17 n857 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_57 n8044 CLK \AES_Comp_ENCa/KrgX_57 n910 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_25 n8076 CLK \AES_Comp_ENCa/KrgX_25 n876 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_33 n8068 CLK \AES_Comp_ENCa/KrgX_33 n886 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_42 n8059 CLK \AES_Comp_ENCa/KrgX_42 n895 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_10 n8091 CLK \AES_Comp_ENCa/KrgX_10 n841 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_51 n8050 CLK \AES_Comp_ENCa/KrgX_51 n904 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_19 n8082 CLK \AES_Comp_ENCa/KrgX_19 n861 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_59 n8042 CLK \AES_Comp_ENCa/KrgX_59 n912 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_27 n8074 CLK \AES_Comp_ENCa/KrgX_27 n879 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_91 n8010 CLK \AES_Comp_ENCa/KrgX_91 n944 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_123 n7978 CLK \AES_Comp_ENCa/KrgX_123 n976 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_60 n8041 CLK \AES_Comp_ENCa/KrgX_60 n913 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_28 n8073 CLK \AES_Comp_ENCa/KrgX_28 n880 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_35 n8066 CLK \AES_Comp_ENCa/KrgX_35 n888 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_3 n8098 CLK \AES_Comp_ENCa/KrgX_3 n827 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_45 n8056 CLK \AES_Comp_ENCa/KrgX_45 n898 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_13 n8088 CLK \AES_Comp_ENCa/KrgX_13 n845 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_77 n8024 CLK \AES_Comp_ENCa/KrgX_77 n930 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_109 n7992 CLK \AES_Comp_ENCa/KrgX_109 n962 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_43 n8058 CLK \AES_Comp_ENCa/KrgX_43 n896 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_11 n8090 CLK \AES_Comp_ENCa/KrgX_11 n842 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_50 n8051 CLK \AES_Comp_ENCa/KrgX_50 n903 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_18 n8083 CLK \AES_Comp_ENCa/KrgX_18 n860 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_63 n8038 CLK \AES_Comp_ENCa/KrgX_63 n916 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_31 n8070 CLK \AES_Comp_ENCa/KrgX_31 n884 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_37 n8064 CLK \AES_Comp_ENCa/KrgX_37 n890 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_5 n8096 CLK \AES_Comp_ENCa/KrgX_5 n830 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_46 n8055 CLK \AES_Comp_ENCa/KrgX_46 n899 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_14 n8087 CLK \AES_Comp_ENCa/KrgX_14 n846 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_54 n8047 CLK \AES_Comp_ENCa/KrgX_54 n907 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_22 n8079 CLK \AES_Comp_ENCa/KrgX_22 n866 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_58 n8043 CLK \AES_Comp_ENCa/KrgX_58 n911 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_26 n8075 CLK \AES_Comp_ENCa/KrgX_26 n878 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_34 n8067 CLK \AES_Comp_ENCa/KrgX_34 n887 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_2 n8099 CLK \AES_Comp_ENCa/KrgX_2 n826 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_47 n8054 CLK \AES_Comp_ENCa/KrgX_47 n900 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_15 n8086 CLK \AES_Comp_ENCa/KrgX_15 n847 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_53 n8048 CLK \AES_Comp_ENCa/KrgX_53 n906 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_21 n8080 CLK \AES_Comp_ENCa/KrgX_21 n865 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_62 n8039 CLK \AES_Comp_ENCa/KrgX_62 n915 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_30 n8071 CLK \AES_Comp_ENCa/KrgX_30 n883 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_38 n8063 CLK \AES_Comp_ENCa/KrgX_38 n891 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_6 n8095 CLK \AES_Comp_ENCa/KrgX_6 n831 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_44 n8057 CLK \AES_Comp_ENCa/KrgX_44 n897 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_12 n8089 CLK \AES_Comp_ENCa/KrgX_12 n844 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_52 n8049 CLK \AES_Comp_ENCa/KrgX_52 n905 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_20 n8081 CLK \AES_Comp_ENCa/KrgX_20 n864 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_84 n8017 CLK \AES_Comp_ENCa/KrgX_84 n937 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_116 n7985 CLK \AES_Comp_ENCa/KrgX_116 n969 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_55 n8046 CLK \AES_Comp_ENCa/KrgX_55 n908 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_23 n8078 CLK \AES_Comp_ENCa/KrgX_23 n867 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_61 n8040 CLK \AES_Comp_ENCa/KrgX_61 n914 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_29 n8072 CLK \AES_Comp_ENCa/KrgX_29 n882 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_39 n8062 CLK \AES_Comp_ENCa/KrgX_39 n892 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_7 n8094 CLK \AES_Comp_ENCa/KrgX_7 n832 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_71 n8030 CLK \AES_Comp_ENCa/KrgX_71 n924 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_103 n7998 CLK \AES_Comp_ENCa/KrgX_103 n956 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_93 n8008 CLK \AES_Comp_ENCa/KrgX_93 n946 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_125 n7976 CLK \AES_Comp_ENCa/KrgX_125 n978 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_87 n8014 CLK \AES_Comp_ENCa/KrgX_87 n940 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_119 n7982 CLK \AES_Comp_ENCa/KrgX_119 n972 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_76 n8025 CLK \AES_Comp_ENCa/KrgX_76 n929 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_108 n7993 CLK \AES_Comp_ENCa/KrgX_108 n961 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_70 n8031 CLK \AES_Comp_ENCa/KrgX_70 n923 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_102 n7999 CLK \AES_Comp_ENCa/KrgX_102 n955 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_94 n8007 CLK \AES_Comp_ENCa/KrgX_94 n947 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_126 n7975 CLK \AES_Comp_ENCa/KrgX_126 n979 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_85 n8016 CLK \AES_Comp_ENCa/KrgX_85 n938 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_117 n7984 CLK \AES_Comp_ENCa/KrgX_117 n970 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_79 n8022 CLK \AES_Comp_ENCa/KrgX_79 n932 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_111 n7990 CLK \AES_Comp_ENCa/KrgX_111 n964 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_66 n8035 CLK \AES_Comp_ENCa/KrgX_66 n919 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_98 n8003 CLK \AES_Comp_ENCa/KrgX_98 n951 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_90 n8011 CLK \AES_Comp_ENCa/KrgX_90 n943 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_122 n7979 CLK \AES_Comp_ENCa/KrgX_122 n975 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_86 n8015 CLK \AES_Comp_ENCa/KrgX_86 n939 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_118 n7983 CLK \AES_Comp_ENCa/KrgX_118 n971 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_78 n8023 CLK \AES_Comp_ENCa/KrgX_78 n931 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_110 n7991 CLK \AES_Comp_ENCa/KrgX_110 n963 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_69 n8032 CLK \AES_Comp_ENCa/KrgX_69 n922 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_101 n8000 CLK \AES_Comp_ENCa/KrgX_101 n954 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_95 n8006 CLK \AES_Comp_ENCa/KrgX_95 n948 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_127 n7974 CLK \AES_Comp_ENCa/KrgX_127 n980 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_82 n8019 CLK \AES_Comp_ENCa/KrgX_82 n935 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_114 n7987 CLK \AES_Comp_ENCa/KrgX_114 n967 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_75 n8026 CLK \AES_Comp_ENCa/KrgX_75 n928 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_107 n7994 CLK \AES_Comp_ENCa/KrgX_107 n960 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_67 n8034 CLK \AES_Comp_ENCa/KrgX_67 n920 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_99 n8002 CLK \AES_Comp_ENCa/KrgX_99 n952 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_92 n8009 CLK \AES_Comp_ENCa/KrgX_92 n945 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_124 n7977 CLK \AES_Comp_ENCa/KrgX_124 n977 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_83 n8018 CLK \AES_Comp_ENCa/KrgX_83 n936 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_115 n7986 CLK \AES_Comp_ENCa/KrgX_115 n968 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_74 n8027 CLK \AES_Comp_ENCa/KrgX_74 n927 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_106 n7995 CLK \AES_Comp_ENCa/KrgX_106 n959 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_65 n8036 CLK \AES_Comp_ENCa/KrgX_65 n918 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_97 n8004 CLK \AES_Comp_ENCa/KrgX_97 n950 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_89 n8012 CLK \AES_Comp_ENCa/KrgX_89 n942 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_121 n7980 CLK \AES_Comp_ENCa/KrgX_121 n974 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_81 n8020 CLK \AES_Comp_ENCa/KrgX_81 n934 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_113 n7988 CLK \AES_Comp_ENCa/KrgX_113 n966 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_73 n8028 CLK \AES_Comp_ENCa/KrgX_73 n926 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_105 n7996 CLK \AES_Comp_ENCa/KrgX_105 n958 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_68 n8033 CLK \AES_Comp_ENCa/KrgX_68 n921 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_100 n8001 CLK \AES_Comp_ENCa/KrgX_100 n953 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_32 n8069 CLK \AES_Comp_ENCa/KrgX_32 n885 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_64 n8037 CLK \AES_Comp_ENCa/KrgX_64 n917 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_96 n8005 CLK \AES_Comp_ENCa/KrgX_96 n949 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_88 n8013 CLK \AES_Comp_ENCa/KrgX_88 n941 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_120 n7981 CLK \AES_Comp_ENCa/KrgX_120 n973 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_80 n8021 CLK \AES_Comp_ENCa/KrgX_80 n933 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_112 n7989 CLK \AES_Comp_ENCa/KrgX_112 n965 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_72 n8029 CLK \AES_Comp_ENCa/KrgX_72 n925 VDD GND DFF_X1
xAES_Comp_ENCa/KrgX_reg_104 n7997 CLK \AES_Comp_ENCa/KrgX_104 n957 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_0 n7973 CLK Dout_E_0 n188 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_97 n7876 CLK Dout_E_97 n593 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_64 n7909 CLK Dout_E_64 n483 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_35 n7938 CLK Dout_E_35 n390 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_3 n7970 CLK Dout_E_3 n192 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_107 n7866 CLK Dout_E_107 n622 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_43 n7930 CLK Dout_E_43 n413 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_117 n7856 CLK Dout_E_117 n654 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_16 n7957 CLK Dout_E_16 n301 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_51 n7922 CLK Dout_E_51 n437 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_80 n7893 CLK Dout_E_80 n538 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_115 n7858 CLK Dout_E_115 n651 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_17 n7956 CLK Dout_E_17 n303 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_48 n7925 CLK Dout_E_48 n433 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_81 n7892 CLK Dout_E_81 n539 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_112 n7861 CLK Dout_E_112 n643 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_19 n7954 CLK Dout_E_19 n307 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_49 n7924 CLK Dout_E_49 n434 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_89 n7884 CLK Dout_E_89 n563 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_92 n7881 CLK Dout_E_92 n568 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_91 n7882 CLK Dout_E_91 n566 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_66 n7907 CLK Dout_E_66 n489 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_32 n7941 CLK Dout_E_32 n386 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_7 n7966 CLK Dout_E_7 n197 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_127 n7846 CLK Dout_E_127 n680 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_96 n7877 CLK Dout_E_96 n591 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_68 n7905 CLK Dout_E_68 n492 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_59 n7914 CLK Dout_E_59 n463 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_41 n7932 CLK Dout_E_41 n411 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_104 n7869 CLK Dout_E_104 n617 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_45 n7928 CLK Dout_E_45 n416 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_105 n7868 CLK Dout_E_105 n618 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_58 n7915 CLK Dout_E_58 n462 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_42 n7931 CLK Dout_E_42 n412 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_106 n7867 CLK Dout_E_106 n621 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_40 n7933 CLK Dout_E_40 n409 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_108 n7865 CLK Dout_E_108 n625 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_33 n7940 CLK Dout_E_33 n388 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_31 n7942 CLK Dout_E_31 n369 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_25 n7948 CLK Dout_E_25 n362 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_1 n7972 CLK Dout_E_1 n190 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_100 n7873 CLK Dout_E_100 n597 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_88 n7885 CLK Dout_E_88 n561 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_70 n7903 CLK Dout_E_70 n494 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_34 n7939 CLK Dout_E_34 n389 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_2 n7971 CLK Dout_E_2 n191 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_98 n7875 CLK Dout_E_98 n594 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_75 n7898 CLK Dout_E_75 n516 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_11 n7962 CLK Dout_E_11 n249 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_85 n7888 CLK Dout_E_85 n544 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_120 n7853 CLK Dout_E_120 n668 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_122 n7851 CLK Dout_E_122 n673 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_103 n7870 CLK Dout_E_103 n600 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_65 n7908 CLK Dout_E_65 n485 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_36 n7937 CLK Dout_E_36 n392 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_18 n7955 CLK Dout_E_18 n306 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_62 n7911 CLK Dout_E_62 n467 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_60 n7913 CLK Dout_E_60 n465 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_37 n7936 CLK Dout_E_37 n393 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_24 n7949 CLK Dout_E_24 n361 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_27 n7946 CLK Dout_E_27 n365 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_28 n7945 CLK Dout_E_28 n366 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_26 n7947 CLK Dout_E_26 n364 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_4 n7969 CLK Dout_E_4 n194 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_102 n7871 CLK Dout_E_102 n599 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_90 n7883 CLK Dout_E_90 n565 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_72 n7901 CLK Dout_E_72 n511 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_9 n7964 CLK Dout_E_9 n245 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_76 n7897 CLK Dout_E_76 n517 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_13 n7960 CLK Dout_E_13 n253 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_73 n7900 CLK Dout_E_73 n513 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_8 n7965 CLK Dout_E_8 n243 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_74 n7899 CLK Dout_E_74 n515 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_14 n7959 CLK Dout_E_14 n254 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_77 n7896 CLK Dout_E_77 n518 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_12 n7961 CLK Dout_E_12 n252 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_83 n7890 CLK Dout_E_83 n542 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_113 n7860 CLK Dout_E_113 n647 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_21 n7952 CLK Dout_E_21 n310 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_50 n7923 CLK Dout_E_50 n436 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_82 n7891 CLK Dout_E_82 n541 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_114 n7859 CLK Dout_E_114 n650 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_6 n7967 CLK Dout_E_6 n196 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_99 n7874 CLK Dout_E_99 n595 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_87 n7886 CLK Dout_E_87 n546 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_116 n7857 CLK dummy7 n653 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_15 n7958 CLK Dout_E_15 n255 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_84 n7889 CLK Dout_E_84 n543 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_126 n7847 CLK Dout_E_126 n679 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_121 n7852 CLK Dout_E_121 n669 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_123 n7850 CLK Dout_E_123 n674 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_111 n7862 CLK Dout_E_111 n628 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_44 n7929 CLK Dout_E_44 n415 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_119 n7854 CLK Dout_E_119 n656 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_10 n7963 CLK Dout_E_10 n248 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_94 n7879 CLK Dout_E_94 n571 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_67 n7906 CLK Dout_E_67 n490 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_39 n7934 CLK Dout_E_39 n395 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_30 n7943 CLK Dout_E_30 n368 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_5 n7968 CLK Dout_E_5 n195 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_118 n7855 CLK Dout_E_118 n655 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_20 n7953 CLK Dout_E_20 n309 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_52 n7921 CLK Dout_E_52 n440 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_93 n7880 CLK Dout_E_93 n570 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_69 n7904 CLK Dout_E_69 n493 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_38 n7935 CLK Dout_E_38 n394 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_29 n7944 CLK Dout_E_29 n367 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_22 n7951 CLK Dout_E_22 n311 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_53 n7920 CLK Dout_E_53 n441 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_71 n7902 CLK Dout_E_71 n495 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_61 n7912 CLK Dout_E_61 n466 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_57 n7916 CLK Dout_E_57 n460 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_56 n7917 CLK Dout_E_56 n459 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_47 n7926 CLK Dout_E_47 n418 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_109 n7864 CLK Dout_E_109 n626 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_54 n7919 CLK Dout_E_54 n442 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_79 n7894 CLK Dout_E_79 n520 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_23 n7950 CLK Dout_E_23 n312 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_63 n7910 CLK Dout_E_63 n468 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_46 n7927 CLK Dout_E_46 n417 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_55 n7918 CLK Dout_E_55 n443 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_95 n7878 CLK Dout_E_95 n572 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_86 n7887 CLK Dout_E_86 n545 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_124 n7849 CLK Dout_E_124 n677 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_125 n7848 CLK Dout_E_125 n678 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_110 n7863 CLK Dout_E_110 n627 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_101 n7872 CLK Dout_E_101 n598 VDD GND DFF_X1
xAES_Comp_ENCa/Drg_reg_78 n7895 CLK Dout_E_78 n519 VDD GND DFF_X1
xAES_Comp_ENCa/Dvldrg_reg n8111 CLK Dvld_E n809 VDD GND DFF_X1
xDvld_reg_reg n8110 CLK Dvld_reg dummy8 VDD GND DFF_X1
xU4692 n996 n997 n992 VDD GND XOR2_X1
xU4693 n998 n999 n997 VDD GND XOR2_X1
xU4694 n1000 n1001 n999 VDD GND XOR2_X1
xU4695 n1002 n1003 n996 VDD GND XOR2_X1
xU4696 n1004 n153 n1003 VDD GND XOR2_X1
xU4697 n808 Din_127 n1008 VDD GND XOR2_X1
xU4698 n1022 n1023 n1017 VDD GND XOR2_X1
xU4699 n661 n1024 n1023 VDD GND XOR2_X1
xU4700 n1025 n1026 n1024 VDD GND XOR2_X1
xU4701 n1027 n998 n1022 VDD GND XOR2_X1
xU4702 n532 n1028 n998 VDD GND XOR2_X1
xU4703 n1029 n405 n1027 VDD GND XOR2_X1
xU4704 n807 Din_126 n1032 VDD GND XOR2_X1
xU4705 n1045 n1046 n1041 VDD GND XOR2_X1
xU4706 n398 n1047 n1046 VDD GND XOR2_X1
xU4707 n522 n1048 n1047 VDD GND XOR2_X1
xU4708 n161 n1049 n1045 VDD GND XOR2_X1
xU4709 n1050 n662 n1049 VDD GND XOR2_X1
xU4710 n806 Din_125 n1053 VDD GND XOR2_X1
xU4711 n1066 n1067 n1062 VDD GND XOR2_X1
xU4712 n1068 n1069 n1067 VDD GND XOR2_X1
xU4713 n1070 n1071 n1069 VDD GND XOR2_X1
xU4714 n1072 n1073 n1068 VDD GND XOR2_X1
xU4715 n1074 n1075 n1066 VDD GND XOR2_X1
xU4716 n1050 n1076 n1075 VDD GND XOR2_X1
xU4717 n1077 n1078 n1074 VDD GND XOR2_X1
xU4718 n805 Din_124 n1081 VDD GND XOR2_X1
xU4719 n1094 n1095 n1090 VDD GND XOR2_X1
xU4720 n1096 n1097 n1095 VDD GND XOR2_X1
xU4721 n1098 n1099 n1097 VDD GND XOR2_X1
xU4722 n1100 n1101 n1094 VDD GND XOR2_X1
xU4723 n1102 n1103 n1101 VDD GND XOR2_X1
xU4724 n804 Din_123 n1106 VDD GND XOR2_X1
xU4725 n1119 n1120 n1115 VDD GND XOR2_X1
xU4726 n1121 n1122 n1120 VDD GND XOR2_X1
xU4727 n1123 n1124 n1122 VDD GND XOR2_X1
xU4728 n660 n1125 n1121 VDD GND XOR2_X1
xU4729 n1126 n1127 n1119 VDD GND XOR2_X1
xU4730 n1001 n1128 n1127 VDD GND XOR2_X1
xU4731 n1129 n1103 n1001 VDD GND XOR2_X1
xU4732 n1130 n1131 n1126 VDD GND XOR2_X1
xU4733 n803 Din_122 n1134 VDD GND XOR2_X1
xU4734 n1147 n1148 n1142 VDD GND XOR2_X1
xU4735 n1149 n1150 n1148 VDD GND XOR2_X1
xU4736 n1098 n1151 n1150 VDD GND XOR2_X1
xU4737 n1152 n1153 n1098 VDD GND XOR2_X1
xU4738 n1154 n1155 n1147 VDD GND XOR2_X1
xU4739 n802 Din_121 n1158 VDD GND XOR2_X1
xU4740 n1171 n1172 n1167 VDD GND XOR2_X1
xU4741 n396 n171 n1172 VDD GND XOR2_X1
xU4742 n1173 n1174 n1171 VDD GND XOR2_X1
xU4743 n1175 n533 n1174 VDD GND XOR2_X1
xU4744 n801 Din_120 n1178 VDD GND XOR2_X1
xU4745 n1191 n1004 n1186 VDD GND XOR2_X1
xU4746 n1192 n1193 n1187 VDD GND XOR2_X1
xU4747 n990 n1194 n1193 VDD GND XOR2_X1
xU4748 n1195 n153 n1194 VDD GND XOR2_X1
xU4749 n1197 n1175 n990 VDD GND XOR2_X1
xU4750 n1198 n1199 n1192 VDD GND XOR2_X1
xU4751 n1200 n1201 n1199 VDD GND XOR2_X1
xU4752 n800 Din_119 n1204 VDD GND XOR2_X1
xU4753 n1029 n1216 n1201 VDD GND XOR2_X1
xU4754 n1217 n1218 n1212 VDD GND XOR2_X1
xU4755 n1026 n1219 n1218 VDD GND XOR2_X1
xU4756 n1128 n1195 n1219 VDD GND XOR2_X1
xU4757 n1220 n1221 n1026 VDD GND XOR2_X1
xU4758 n523 n1222 n1217 VDD GND XOR2_X1
xU4759 n663 n1223 n1222 VDD GND XOR2_X1
xU4760 n1224 n1225 n1021 VDD GND XOR2_X1
xU4761 n799 Din_118 n1228 VDD GND XOR2_X1
xU4762 n1241 n1242 n1236 VDD GND XOR2_X1
xU4763 n161 n1243 n1242 VDD GND XOR2_X1
xU4764 n661 n1244 n1243 VDD GND XOR2_X1
xU4765 n528 n1245 n1241 VDD GND XOR2_X1
xU4766 n1246 n397 n1245 VDD GND XOR2_X1
xU4767 n798 Din_117 n1249 VDD GND XOR2_X1
xU4768 n1262 n1263 n1258 VDD GND XOR2_X1
xU4769 n1264 n1265 n1263 VDD GND XOR2_X1
xU4770 n166 n1266 n1265 VDD GND XOR2_X1
xU4771 n1061 n1244 n1264 VDD GND XOR2_X1
xU4772 n1267 n1268 n1262 VDD GND XOR2_X1
xU4773 n1269 n1270 n1268 VDD GND XOR2_X1
xU4774 n1271 n1272 n1267 VDD GND XOR2_X1
xU4775 n797 Din_116 n1275 VDD GND XOR2_X1
xU4776 n1288 n1289 n1284 VDD GND XOR2_X1
xU4777 n1290 n1291 n1289 VDD GND XOR2_X1
xU4778 n1292 n1293 n1291 VDD GND XOR2_X1
xU4779 n1294 n1099 n1290 VDD GND XOR2_X1
xU4780 n179 n1130 n1099 VDD GND XOR2_X1
xU4781 n1295 n1296 n1288 VDD GND XOR2_X1
xU4782 n1297 n1298 n1296 VDD GND XOR2_X1
xU4783 n1029 n1299 n1295 VDD GND XOR2_X1
xU4784 n796 Din_115 n1302 VDD GND XOR2_X1
xU4785 n1125 n1315 n1310 VDD GND XOR2_X1
xU4786 n1029 n1004 n1125 VDD GND XOR2_X1
xU4787 n1316 n1317 n1311 VDD GND XOR2_X1
xU4788 n1318 n1319 n1317 VDD GND XOR2_X1
xU4789 n1198 n1114 n1319 VDD GND XOR2_X1
xU4790 n1320 n1321 n1114 VDD GND XOR2_X1
xU4791 n1197 n1322 n1321 VDD GND XOR2_X1
xU4792 n148 n1297 n1198 VDD GND XOR2_X1
xU4793 n1123 n1323 n1316 VDD GND XOR2_X1
xU4794 n1324 n181 n1323 VDD GND XOR2_X1
xU4795 n795 Din_114 n1327 VDD GND XOR2_X1
xU4796 n1340 n1341 n1336 VDD GND XOR2_X1
xU4797 n1342 n1343 n1341 VDD GND XOR2_X1
xU4798 n660 n1294 n1343 VDD GND XOR2_X1
xU4799 n1270 n1344 n1340 VDD GND XOR2_X1
xU4800 n1173 n1345 n1344 VDD GND XOR2_X1
xU4801 n1346 n1347 n1173 VDD GND XOR2_X1
xU4802 n1348 n1272 n1347 VDD GND XOR2_X1
xU4803 n529 n1153 n1272 VDD GND XOR2_X1
xU4804 n1349 n1350 n1346 VDD GND XOR2_X1
xU4805 n1351 n1050 n1350 VDD GND XOR2_X1
xU4806 n794 Din_113 n1354 VDD GND XOR2_X1
xU4807 n1367 n1368 n1363 VDD GND XOR2_X1
xU4808 n525 n1369 n1368 VDD GND XOR2_X1
xU4809 n1166 n171 n1369 VDD GND XOR2_X1
xU4810 n1270 n1370 n1367 VDD GND XOR2_X1
xU4811 n406 n1004 n1270 VDD GND XOR2_X1
xU4812 n793 Din_112 n1373 VDD GND XOR2_X1
xU4813 n1000 n406 n1381 VDD GND XOR2_X1
xU4814 n1386 n1387 n1382 VDD GND XOR2_X1
xU4815 n1388 n1389 n1387 VDD GND XOR2_X1
xU4816 n1191 n1390 n1389 VDD GND XOR2_X1
xU4817 n1391 n1392 n1386 VDD GND XOR2_X1
xU4818 n1175 n181 n1392 VDD GND XOR2_X1
xU4819 n1076 n1393 n1175 VDD GND XOR2_X1
xU4820 n405 n1394 n1391 VDD GND XOR2_X1
xU4821 n792 Din_111 n1397 VDD GND XOR2_X1
xU4822 n1410 n1411 n1406 VDD GND XOR2_X1
xU4823 n1388 n1412 n1411 VDD GND XOR2_X1
xU4824 n398 n1413 n1412 VDD GND XOR2_X1
xU4825 n1414 n1415 n1388 VDD GND XOR2_X1
xU4826 n1416 n1417 n1410 VDD GND XOR2_X1
xU4827 n1216 n1002 n1417 VDD GND XOR2_X1
xU4828 n1102 n1225 n1002 VDD GND XOR2_X1
xU4829 n791 Din_110 n1420 VDD GND XOR2_X1
xU4830 n1433 n1434 n1429 VDD GND XOR2_X1
xU4831 n1435 n1436 n1434 VDD GND XOR2_X1
xU4832 n661 n1437 n1436 VDD GND XOR2_X1
xU4833 n1076 n1438 n1040 VDD GND XOR2_X1
xU4834 n523 n1439 n1433 VDD GND XOR2_X1
xU4835 n402 n179 n1439 VDD GND XOR2_X1
xU4836 n790 Din_109 n1442 VDD GND XOR2_X1
xU4837 n1454 n1455 n1450 VDD GND XOR2_X1
xU4838 n1456 n1457 n1455 VDD GND XOR2_X1
xU4839 n1257 n1155 n1457 VDD GND XOR2_X1
xU4840 n1294 n1458 n1456 VDD GND XOR2_X1
xU4841 n1459 n1460 n1454 VDD GND XOR2_X1
xU4842 n1061 n1461 n1460 VDD GND XOR2_X1
xU4843 n1462 n1463 n1061 VDD GND XOR2_X1
xU4844 n1464 n1465 n1463 VDD GND XOR2_X1
xU4845 n1466 n1467 n1462 VDD GND XOR2_X1
xU4846 n1468 n1469 n1466 VDD GND XOR2_X1
xU4847 n148 n1437 n1459 VDD GND XOR2_X1
xU4848 n789 Din_108 n1472 VDD GND XOR2_X1
xU4849 n1485 n1486 n1481 VDD GND XOR2_X1
xU4850 n1487 n1488 n1486 VDD GND XOR2_X1
xU4851 n1293 n1124 n1488 VDD GND XOR2_X1
xU4852 n181 n1489 n1124 VDD GND XOR2_X1
xU4853 n1298 n1416 n1220 VDD GND XOR2_X1
xU4854 n1089 n1324 n1293 VDD GND XOR2_X1
xU4855 n182 n1490 n1485 VDD GND XOR2_X1
xU4856 n1491 n1492 n1490 VDD GND XOR2_X1
xU4857 n788 Din_107 n1495 VDD GND XOR2_X1
xU4858 n1508 n1509 n1503 VDD GND XOR2_X1
xU4859 n1510 n1299 n1508 VDD GND XOR2_X1
xU4860 n1511 n1512 n1504 VDD GND XOR2_X1
xU4861 n1513 n1514 n1512 VDD GND XOR2_X1
xU4862 n1515 n1516 n1514 VDD GND XOR2_X1
xU4863 n1517 n1518 n1511 VDD GND XOR2_X1
xU4864 n1315 n1390 n1518 VDD GND XOR2_X1
xU4865 n1491 n533 n1390 VDD GND XOR2_X1
xU4866 n1519 n1320 n1517 VDD GND XOR2_X1
xU4867 n1520 n1521 n1320 VDD GND XOR2_X1
xU4868 n787 Din_106 n1524 VDD GND XOR2_X1
xU4869 n1536 n1537 n1532 VDD GND XOR2_X1
xU4870 n1370 n1538 n1537 VDD GND XOR2_X1
xU4871 n1539 n1318 n1538 VDD GND XOR2_X1
xU4872 n524 n1540 n1318 VDD GND XOR2_X1
xU4873 n1541 n1542 n1370 VDD GND XOR2_X1
xU4874 n1543 n1544 n1542 VDD GND XOR2_X1
xU4875 n1294 n1492 n1544 VDD GND XOR2_X1
xU4876 n1545 n1546 n1541 VDD GND XOR2_X1
xU4877 n1195 n1244 n1546 VDD GND XOR2_X1
xU4878 n660 n1547 n1536 VDD GND XOR2_X1
xU4879 n1129 n182 n1547 VDD GND XOR2_X1
xU4880 n1076 n1096 n1146 VDD GND XOR2_X1
xU4881 n1520 n1548 n1096 VDD GND XOR2_X1
xU4882 n1464 n1549 n1076 VDD GND XOR2_X1
xU4883 n786 Din_105 n1552 VDD GND XOR2_X1
xU4884 n1565 n1566 n1561 VDD GND XOR2_X1
xU4885 n1567 n1568 n1566 VDD GND XOR2_X1
xU4886 n1000 n148 n1568 VDD GND XOR2_X1
xU4887 n406 n1394 n1129 VDD GND XOR2_X1
xU4888 n1569 n1570 n1565 VDD GND XOR2_X1
xU4889 n659 n521 n1570 VDD GND XOR2_X1
xU4890 n664 n1571 n1166 VDD GND XOR2_X1
xU4891 n785 Din_104 n1574 VDD GND XOR2_X1
xU4892 n1196 n1394 n1582 VDD GND XOR2_X1
xU4893 n1587 n1588 n1583 VDD GND XOR2_X1
xU4894 n1589 n1590 n1588 VDD GND XOR2_X1
xU4895 n533 n1322 n1590 VDD GND XOR2_X1
xU4896 n1224 n1549 n1322 VDD GND XOR2_X1
xU4897 n1000 n665 n1589 VDD GND XOR2_X1
xU4898 n1297 n1591 n1000 VDD GND XOR2_X1
xU4899 n173 n1592 n1587 VDD GND XOR2_X1
xU4900 n525 n1593 n1592 VDD GND XOR2_X1
xU4901 n1269 n1103 n1191 VDD GND XOR2_X1
xU4902 n784 Din_103 n1596 VDD GND XOR2_X1
xU4903 n1416 n1221 n1604 VDD GND XOR2_X1
xU4904 n1609 n1610 n1605 VDD GND XOR2_X1
xU4905 n1513 n1611 n1610 VDD GND XOR2_X1
xU4906 n1612 n403 n1611 VDD GND XOR2_X1
xU4907 n1298 n405 n1405 VDD GND XOR2_X1
xU4908 n530 n1549 n1513 VDD GND XOR2_X1
xU4909 n1613 n1467 n1549 VDD GND XOR2_X1
xU4910 n1614 n1615 n1467 VDD GND XOR2_X1
xU4911 n1616 n1438 n1609 VDD GND XOR2_X1
xU4912 n1617 n1618 n1438 VDD GND XOR2_X1
xU4913 n1216 n665 n1616 VDD GND XOR2_X1
xU4914 n783 Din_102 n1621 VDD GND XOR2_X1
xU4915 n1633 n1413 n1612 VDD GND XOR2_X1
xU4916 n1634 n1461 n1413 VDD GND XOR2_X1
xU4917 n1635 n1636 n1461 VDD GND XOR2_X1
xU4918 n1637 n1638 n1629 VDD GND XOR2_X1
xU4919 n1428 n1639 n1638 VDD GND XOR2_X1
xU4920 n1613 n1640 n1639 VDD GND XOR2_X1
xU4921 n1223 n1591 n1428 VDD GND XOR2_X1
xU4922 n1641 n1266 n1223 VDD GND XOR2_X1
xU4923 n1642 n1643 n1266 VDD GND XOR2_X1
xU4924 n523 n1644 n1637 VDD GND XOR2_X1
xU4925 n1073 n1089 n1644 VDD GND XOR2_X1
xU4926 n1645 n1521 n1089 VDD GND XOR2_X1
xU4927 n1393 n1548 n1521 VDD GND XOR2_X1
xU4928 n1269 n1025 n1240 VDD GND XOR2_X1
xU4929 n1646 n1077 n1025 VDD GND XOR2_X1
xU4930 n1647 n1648 n1077 VDD GND XOR2_X1
xU4931 n782 Din_101 n1651 VDD GND XOR2_X1
xU4932 n1663 n1664 n1073 VDD GND XOR2_X1
xU4933 n1519 n1458 n1664 VDD GND XOR2_X1
xU4934 n1435 n1665 n1458 VDD GND XOR2_X1
xU4935 n1666 n1667 n1435 VDD GND XOR2_X1
xU4936 n1668 n1669 n1667 VDD GND XOR2_X1
xU4937 Dout_E_1 n1672 n1670 VDD GND XOR2_X1
xU4938 n1673 n184 n1663 VDD GND XOR2_X1
xU4939 n1674 n1675 n1673 VDD GND XOR2_X1
xU4940 n1676 n1677 n1659 VDD GND XOR2_X1
xU4941 n1678 n1679 n1677 VDD GND XOR2_X1
xU4942 n1072 n1465 n1679 VDD GND XOR2_X1
xU4943 n1640 n1680 n1465 VDD GND XOR2_X1
xU4944 n1681 n1682 n1640 VDD GND XOR2_X1
xU4945 n1683 n1684 n1682 VDD GND XOR2_X1
xU4946 n669 n1687 n1685 VDD GND XOR2_X1
xU4947 n1688 n1689 n1072 VDD GND XOR2_X1
xU4948 n1324 n1271 n1689 VDD GND XOR2_X1
xU4949 n1246 n1690 n1271 VDD GND XOR2_X1
xU4950 n1691 n1692 n1246 VDD GND XOR2_X1
xU4951 n1693 n1694 n1692 VDD GND XOR2_X1
xU4952 Dout_E_41 n1697 n1695 VDD GND XOR2_X1
xU4953 n1698 n1699 n1688 VDD GND XOR2_X1
xU4954 n1700 n1701 n1698 VDD GND XOR2_X1
xU4955 n1613 n1618 n1678 VDD GND XOR2_X1
xU4956 n1702 n1703 n1618 VDD GND XOR2_X1
xU4957 n1704 n1705 n1676 VDD GND XOR2_X1
xU4958 n182 n158 n1705 VDD GND XOR2_X1
xU4959 n528 n1706 n1704 VDD GND XOR2_X1
xU4960 n1707 n1708 n1257 VDD GND XOR2_X1
xU4961 n1078 n1130 n1708 VDD GND XOR2_X1
xU4962 n1048 n1709 n1078 VDD GND XOR2_X1
xU4963 n1710 n1711 n1048 VDD GND XOR2_X1
xU4964 n1712 n1713 n1711 VDD GND XOR2_X1
xU4965 n539 n540 n1714 VDD GND XOR2_X1
xU4966 n1716 n1717 n1707 VDD GND XOR2_X1
xU4967 n1718 n1719 n1716 VDD GND XOR2_X1
xU4968 n781 Din_100 n1722 VDD GND XOR2_X1
xU4969 n1735 n1736 n1730 VDD GND XOR2_X1
xU4970 n1737 n1738 n1736 VDD GND XOR2_X1
xU4971 n1100 n1487 n1738 VDD GND XOR2_X1
xU4972 n522 n1519 n1487 VDD GND XOR2_X1
xU4973 n397 n1464 n1100 VDD GND XOR2_X1
xU4974 n1739 n1740 n1735 VDD GND XOR2_X1
xU4975 n1393 n1416 n1740 VDD GND XOR2_X1
xU4976 n1224 n1540 n1739 VDD GND XOR2_X1
xU4977 n780 Din_99 n1743 VDD GND XOR2_X1
xU4978 n1516 n1756 n1751 VDD GND XOR2_X1
xU4979 n1540 n1123 n1756 VDD GND XOR2_X1
xU4980 n1415 n1757 n1123 VDD GND XOR2_X1
xU4981 n1416 n1394 n1516 VDD GND XOR2_X1
xU4982 n1758 n1759 n1416 VDD GND XOR2_X1
xU4983 n1760 n1668 n1759 VDD GND XOR2_X1
xU4984 n190 n1763 n1761 VDD GND XOR2_X1
xU4985 n1766 n1767 n1752 VDD GND XOR2_X1
xU4986 n1149 n1768 n1767 VDD GND XOR2_X1
xU4987 n530 n1464 n1768 VDD GND XOR2_X1
xU4988 n1225 n665 n1464 VDD GND XOR2_X1
xU4989 n1029 n1224 n1102 VDD GND XOR2_X1
xU4990 n1770 n1771 n1224 VDD GND XOR2_X1
xU4991 n1772 n1683 n1771 VDD GND XOR2_X1
xU4992 Dout_E_121 n670 n1773 VDD GND XOR2_X1
xU4993 n1712 n1777 n1029 VDD GND XOR2_X1
xU4994 n1778 n1779 n1777 VDD GND XOR2_X1
xU4995 Dout_E_81 n1784 n1782 VDD GND XOR2_X1
xU4996 n1070 n1342 n1149 VDD GND XOR2_X1
xU4997 n1489 n158 n1342 VDD GND XOR2_X1
xU4998 n1299 n1540 n1489 VDD GND XOR2_X1
xU4999 n1004 n1197 n1070 VDD GND XOR2_X1
xU5000 n1593 n1788 n1766 VDD GND XOR2_X1
xU5001 n1315 n1509 n1788 VDD GND XOR2_X1
xU5002 n1131 n1200 n1509 VDD GND XOR2_X1
xU5003 n1128 n1298 n1200 VDD GND XOR2_X1
xU5004 n1693 n1789 n1298 VDD GND XOR2_X1
xU5005 n1790 n1791 n1789 VDD GND XOR2_X1
xU5006 Dout_E_41 n1796 n1794 VDD GND XOR2_X1
xU5007 n1797 n1798 n1315 VDD GND XOR2_X1
xU5008 n1152 n1028 n1798 VDD GND XOR2_X1
xU5009 n1393 n406 n1593 VDD GND XOR2_X1
xU5010 n1617 n1680 n1393 VDD GND XOR2_X1
xU5011 n779 Din_98 n1807 VDD GND XOR2_X1
xU5012 n1540 n1785 n1815 VDD GND XOR2_X1
xU5013 n1633 n1567 n1785 VDD GND XOR2_X1
xU5014 n1821 n1822 n1816 VDD GND XOR2_X1
xU5015 n1515 n1823 n1822 VDD GND XOR2_X1
xU5016 n1335 n1571 n1823 VDD GND XOR2_X1
xU5017 n1824 n1825 n1571 VDD GND XOR2_X1
xU5018 n1225 n1615 n1824 VDD GND XOR2_X1
xU5019 n1826 n1827 n1801 VDD GND XOR2_X1
xU5020 n1269 n1292 n1335 VDD GND XOR2_X1
xU5021 n1152 n529 n1292 VDD GND XOR2_X1
xU5022 n1130 n1028 n1269 VDD GND XOR2_X1
xU5023 n1050 n1717 n1028 VDD GND XOR2_X1
xU5024 n1349 n1831 n1717 VDD GND XOR2_X1
xU5025 Dout_E_81 n1836 n1834 VDD GND XOR2_X1
xU5026 n1216 n532 n1130 VDD GND XOR2_X1
xU5027 n1155 n1299 n1515 VDD GND XOR2_X1
xU5028 n1492 n1591 n1155 VDD GND XOR2_X1
xU5029 n1128 n1324 n1591 VDD GND XOR2_X1
xU5030 n405 n1195 n1324 VDD GND XOR2_X1
xU5031 n1244 n1699 n1128 VDD GND XOR2_X1
xU5032 n1545 n1843 n1699 VDD GND XOR2_X1
xU5033 Dout_E_41 n1848 n1846 VDD GND XOR2_X1
xU5034 n1737 n1849 n1821 VDD GND XOR2_X1
xU5035 n1569 n1706 n1849 VDD GND XOR2_X1
xU5036 n1850 n1851 n1569 VDD GND XOR2_X1
xU5037 n1852 n1853 n1851 VDD GND XOR2_X1
xU5038 n1854 n1855 n1850 VDD GND XOR2_X1
xU5039 n1414 n1437 n1855 VDD GND XOR2_X1
xU5040 n1567 n1856 n1737 VDD GND XOR2_X1
xU5041 n1520 n1645 n1856 VDD GND XOR2_X1
xU5042 n778 Din_97 n1862 VDD GND XOR2_X1
xU5043 n179 n1539 n1870 VDD GND XOR2_X1
xU5044 n1875 n1853 n1539 VDD GND XOR2_X1
xU5045 n1758 n1666 n1853 VDD GND XOR2_X1
xU5046 n1221 n1880 n1875 VDD GND XOR2_X1
xU5047 n182 n1757 n1734 VDD GND XOR2_X1
xU5048 n1491 n1567 n1757 VDD GND XOR2_X1
xU5049 n1636 n1675 n1567 VDD GND XOR2_X1
xU5050 n1635 n1674 n1852 VDD GND XOR2_X1
xU5051 n1885 n1886 n1871 VDD GND XOR2_X1
xU5052 n396 n1887 n1886 VDD GND XOR2_X1
xU5053 n1196 n1154 n1887 VDD GND XOR2_X1
xU5054 n1888 n1889 n1154 VDD GND XOR2_X1
xU5055 n1071 n1825 n1889 VDD GND XOR2_X1
xU5056 n1770 n1681 n1825 VDD GND XOR2_X1
xU5057 n1775 n1890 n1803 VDD GND XOR2_X1
xU5058 n1548 n1645 n1071 VDD GND XOR2_X1
xU5059 n1702 n1468 n1645 VDD GND XOR2_X1
xU5060 n1703 n1469 n1548 VDD GND XOR2_X1
xU5061 n1614 n1898 n1888 VDD GND XOR2_X1
xU5062 n1769 n1613 n1898 VDD GND XOR2_X1
xU5063 n1900 n1827 n1896 VDD GND XOR2_X1
xU5064 Dout_E_121 n1891 n1899 VDD GND XOR2_X1
xU5065 n1826 n1900 n1890 VDD GND XOR2_X1
xU5066 n1902 n1903 n1894 VDD GND XOR2_X1
xU5067 n1900 n1893 n1903 VDD GND XOR2_X1
xU5068 n1906 n1907 n1904 VDD GND XOR2_X1
xU5069 n1908 n1909 n1907 VDD GND XOR2_X1
xU5070 n1633 n1491 n1196 VDD GND XOR2_X1
xU5071 n1634 n1665 n1491 VDD GND XOR2_X1
xU5072 n1764 n1876 n1878 VDD GND XOR2_X1
xU5073 n1519 n1415 n1633 VDD GND XOR2_X1
xU5074 n1437 n184 n1415 VDD GND XOR2_X1
xU5075 n1854 n1880 n1914 VDD GND XOR2_X1
xU5076 n1762 n185 n1883 VDD GND XOR2_X1
xU5077 n1922 n1923 n1921 VDD GND XOR2_X1
xU5078 Dout_E_1 n1877 n1920 VDD GND XOR2_X1
xU5079 n1221 n1414 n1519 VDD GND XOR2_X1
xU5080 n1922 n1925 n1876 VDD GND XOR2_X1
xU5081 n1927 n1928 n1918 VDD GND XOR2_X1
xU5082 n1929 n1930 n1928 VDD GND XOR2_X1
xU5083 n397 n1345 n1560 VDD GND XOR2_X1
xU5084 n1932 n1543 n1345 VDD GND XOR2_X1
xU5085 n404 n1691 n1543 VDD GND XOR2_X1
xU5086 n1842 n1843 n1932 VDD GND XOR2_X1
xU5087 n1696 n1935 n1799 VDD GND XOR2_X1
xU5088 n1294 n1131 n1480 VDD GND XOR2_X1
xU5089 n1297 n1492 n1131 VDD GND XOR2_X1
xU5090 n1643 n1701 n1492 VDD GND XOR2_X1
xU5091 n1641 n1690 n1297 VDD GND XOR2_X1
xU5092 n1940 n1941 n1935 VDD GND XOR2_X1
xU5093 n1792 n1840 n1933 VDD GND XOR2_X1
xU5094 n1943 n1940 n1840 VDD GND XOR2_X1
xU5095 n1642 n1700 n1294 VDD GND XOR2_X1
xU5096 n1949 n1950 n1944 VDD GND XOR2_X1
xU5097 n1951 n1952 n1950 VDD GND XOR2_X1
xU5098 n1795 n1847 n1844 VDD GND XOR2_X1
xU5099 n1943 n1941 n1847 VDD GND XOR2_X1
xU5100 n407 n1958 n1949 VDD GND XOR2_X1
xU5101 n408 n1796 n1958 VDD GND XOR2_X1
xU5102 n1960 n1961 n1954 VDD GND XOR2_X1
xU5103 n1951 n1962 n1961 VDD GND XOR2_X1
xU5104 n1964 n1965 n1957 VDD GND XOR2_X1
xU5105 n1845 n1966 n1965 VDD GND XOR2_X1
xU5106 n1967 n1968 n1964 VDD GND XOR2_X1
xU5107 n1969 n1970 n1963 VDD GND XOR2_X1
xU5108 n1968 n1971 n1969 VDD GND XOR2_X1
xU5109 n1966 n1972 n1960 VDD GND XOR2_X1
xU5110 n1934 n1970 n1972 VDD GND XOR2_X1
xU5111 n1973 n1974 n1970 VDD GND XOR2_X1
xU5112 n1975 n1976 n1966 VDD GND XOR2_X1
xU5113 n1948 n1977 n1956 VDD GND XOR2_X1
xU5114 n1962 n1952 n1977 VDD GND XOR2_X1
xU5115 n1971 n1979 n1955 VDD GND XOR2_X1
xU5116 n1980 n1959 n1979 VDD GND XOR2_X1
xU5117 n1975 n1981 n1959 VDD GND XOR2_X1
xU5118 Dout_E_40 n1796 n1982 VDD GND XOR2_X1
xU5119 n1697 n1967 n1971 VDD GND XOR2_X1
xU5120 n1845 n1934 n1697 VDD GND XOR2_X1
xU5121 n410 n1983 n1978 VDD GND XOR2_X1
xU5122 n1793 n408 n1983 VDD GND XOR2_X1
xU5123 n1985 n1974 n1984 VDD GND XOR2_X1
xU5124 Dout_E_40 n1987 n1986 VDD GND XOR2_X1
xU5125 Dout_E_46 n1953 n1938 VDD GND XOR2_X1
xU5126 Dout_E_40 n1848 n1953 VDD GND XOR2_X1
xU5127 Dout_E_45 n1988 n1848 VDD GND XOR2_X1
xU5128 Dout_E_45 Dout_E_47 n1793 VDD GND XOR2_X1
xU5129 n1980 n1967 n1989 VDD GND XOR2_X1
xU5130 Dout_E_43 n414 n1990 VDD GND XOR2_X1
xU5131 Dout_E_41 n1991 n1839 VDD GND XOR2_X1
xU5132 n1993 n1994 n1945 VDD GND XOR2_X1
xU5133 n1934 n1995 n1993 VDD GND XOR2_X1
xU5134 n1996 n1997 n1992 VDD GND XOR2_X1
xU5135 n1994 n1796 n1997 VDD GND XOR2_X1
xU5136 n414 n1988 n1796 VDD GND XOR2_X1
xU5137 n1968 n1980 n1994 VDD GND XOR2_X1
xU5138 n1987 n1999 n1998 VDD GND XOR2_X1
xU5139 Dout_E_47 Dout_E_42 n1999 VDD GND XOR2_X1
xU5140 n1991 n1987 n1946 VDD GND XOR2_X1
xU5141 n417 n411 n1987 VDD GND XOR2_X1
xU5142 Dout_E_44 n2001 n2000 VDD GND XOR2_X1
xU5143 n2002 n2003 n1948 VDD GND XOR2_X1
xU5144 n2004 n1996 n2003 VDD GND XOR2_X1
xU5145 n1973 n1985 n1996 VDD GND XOR2_X1
xU5146 Dout_E_41 n2005 n1939 VDD GND XOR2_X1
xU5147 n1845 n2001 n1841 VDD GND XOR2_X1
xU5148 Dout_E_41 n1988 n2001 VDD GND XOR2_X1
xU5149 Dout_E_47 n1934 n1988 VDD GND XOR2_X1
xU5150 Dout_E_42 Dout_E_43 n1934 VDD GND XOR2_X1
xU5151 Dout_E_45 n414 n1845 VDD GND XOR2_X1
xU5152 n415 Dout_E_46 n2004 VDD GND XOR2_X1
xU5153 n418 n1995 n2002 VDD GND XOR2_X1
xU5154 n1981 n1976 n1995 VDD GND XOR2_X1
xU5155 Dout_E_43 n2009 n1942 VDD GND XOR2_X1
xU5156 Dout_E_42 n2009 n2008 VDD GND XOR2_X1
xU5157 n415 n418 n2009 VDD GND XOR2_X1
xU5158 n2005 n1991 n1800 VDD GND XOR2_X1
xU5159 Dout_E_42 Dout_E_45 n1991 VDD GND XOR2_X1
xU5160 Dout_E_40 Dout_E_44 n2005 VDD GND XOR2_X1
xU5161 Dout_E_40 n2011 n2010 VDD GND XOR2_X1
xU5162 Dout_E_46 Dout_E_43 n2011 VDD GND XOR2_X1
xU5163 n1362 n1706 n1885 VDD GND XOR2_X1
xU5164 n1394 n1197 n1706 VDD GND XOR2_X1
xU5165 n1902 n2013 n1828 VDD GND XOR2_X1
xU5166 n1826 n1859 n2013 VDD GND XOR2_X1
xU5167 n2015 n2016 n1906 VDD GND XOR2_X1
xU5168 n2017 n2018 n2016 VDD GND XOR2_X1
xU5169 n680 n2019 n2015 VDD GND XOR2_X1
xU5170 n2021 n2022 n2014 VDD GND XOR2_X1
xU5171 n2023 n1908 n2022 VDD GND XOR2_X1
xU5172 n1776 n2026 n2024 VDD GND XOR2_X1
xU5173 n2027 n2028 n2026 VDD GND XOR2_X1
xU5174 Dout_E_127 Dout_E_125 n1776 VDD GND XOR2_X1
xU5175 n1827 n1858 n1902 VDD GND XOR2_X1
xU5176 n2028 n2030 n2021 VDD GND XOR2_X1
xU5177 n2031 n2032 n2030 VDD GND XOR2_X1
xU5178 n2033 n2034 n2028 VDD GND XOR2_X1
xU5179 n2027 n2035 n2025 VDD GND XOR2_X1
xU5180 n2032 n1687 n2035 VDD GND XOR2_X1
xU5181 n2036 n2037 n2032 VDD GND XOR2_X1
xU5182 n2038 n2039 n2027 VDD GND XOR2_X1
xU5183 n2040 n1905 n2029 VDD GND XOR2_X1
xU5184 n2041 n2042 n1905 VDD GND XOR2_X1
xU5185 n2043 n2044 n2042 VDD GND XOR2_X1
xU5186 n2047 n2048 n2046 VDD GND XOR2_X1
xU5187 n2044 n2049 n2048 VDD GND XOR2_X1
xU5188 n2036 n2050 n2044 VDD GND XOR2_X1
xU5189 Dout_E_120 n670 n2051 VDD GND XOR2_X1
xU5190 n1891 Dout_E_120 n1895 VDD GND XOR2_X1
xU5191 n1687 n2052 n2045 VDD GND XOR2_X1
xU5192 n2041 n2047 n2052 VDD GND XOR2_X1
xU5193 n2053 n2039 n2047 VDD GND XOR2_X1
xU5194 Dout_E_123 n676 n2054 VDD GND XOR2_X1
xU5195 Dout_E_125 n2055 n1857 VDD GND XOR2_X1
xU5196 n2056 n2033 n2041 VDD GND XOR2_X1
xU5197 Dout_E_121 n2058 n2057 VDD GND XOR2_X1
xU5198 n1891 n2058 n1897 VDD GND XOR2_X1
xU5199 Dout_E_125 n2059 n1891 VDD GND XOR2_X1
xU5200 n2049 n672 n1687 VDD GND XOR2_X1
xU5201 n2017 n2061 n2020 VDD GND XOR2_X1
xU5202 n672 n2062 n2061 VDD GND XOR2_X1
xU5203 n2037 n2050 n2017 VDD GND XOR2_X1
xU5204 Dout_E_122 n2064 n2063 VDD GND XOR2_X1
xU5205 Dout_E_123 n2064 n1804 VDD GND XOR2_X1
xU5206 n677 n680 n2064 VDD GND XOR2_X1
xU5207 n2066 n2067 n2012 VDD GND XOR2_X1
xU5208 n673 n678 n2066 VDD GND XOR2_X1
xU5209 Dout_E_123 n2058 n2065 VDD GND XOR2_X1
xU5210 n668 n679 n2058 VDD GND XOR2_X1
xU5211 n2018 n2068 n2060 VDD GND XOR2_X1
xU5212 n670 n2062 n2068 VDD GND XOR2_X1
xU5213 n2053 n2038 n2062 VDD GND XOR2_X1
xU5214 Dout_E_127 n2070 n2069 VDD GND XOR2_X1
xU5215 Dout_E_125 n2070 n1892 VDD GND XOR2_X1
xU5216 Dout_E_126 n2055 n2070 VDD GND XOR2_X1
xU5217 n673 n669 n2055 VDD GND XOR2_X1
xU5218 Dout_E_124 n2072 n2071 VDD GND XOR2_X1
xU5219 n2019 n2059 n2031 VDD GND XOR2_X1
xU5220 n2056 n2034 n2018 VDD GND XOR2_X1
xU5221 Dout_E_121 n2067 n1802 VDD GND XOR2_X1
xU5222 n668 n677 n2067 VDD GND XOR2_X1
xU5223 n675 n2072 n1901 VDD GND XOR2_X1
xU5224 Dout_E_121 n2059 n2072 VDD GND XOR2_X1
xU5225 n680 n2043 n2059 VDD GND XOR2_X1
xU5226 n673 Dout_E_123 n2043 VDD GND XOR2_X1
xU5227 n678 n676 n2049 VDD GND XOR2_X1
xU5228 n677 Dout_E_126 n2019 VDD GND XOR2_X1
xU5229 n1671 n183 n1931 VDD GND XOR2_X1
xU5230 n1925 n1923 n1915 VDD GND XOR2_X1
xU5231 n1919 n2081 n2076 VDD GND XOR2_X1
xU5232 n2082 n1929 n2081 VDD GND XOR2_X1
xU5233 n2084 n2085 n2079 VDD GND XOR2_X1
xU5234 n1879 n2086 n2084 VDD GND XOR2_X1
xU5235 n187 n2087 n2083 VDD GND XOR2_X1
xU5236 n2085 n1763 n2087 VDD GND XOR2_X1
xU5237 n2088 n2089 n2085 VDD GND XOR2_X1
xU5238 n2091 n2092 n1919 VDD GND XOR2_X1
xU5239 n1879 n2093 n2092 VDD GND XOR2_X1
xU5240 n2080 n2094 n2078 VDD GND XOR2_X1
xU5241 n2082 n1930 n2094 VDD GND XOR2_X1
xU5242 n2096 n2097 n2077 VDD GND XOR2_X1
xU5243 n2089 n2098 n2097 VDD GND XOR2_X1
xU5244 n2099 n2100 n2095 VDD GND XOR2_X1
xU5245 n1765 n186 n2100 VDD GND XOR2_X1
xU5246 Dout_E_7 Dout_E_5 n1765 VDD GND XOR2_X1
xU5247 n2101 n2089 n2099 VDD GND XOR2_X1
xU5248 Dout_E_7 n2103 n2102 VDD GND XOR2_X1
xU5249 Dout_E_5 n2103 n1882 VDD GND XOR2_X1
xU5250 Dout_E_6 n2104 n2103 VDD GND XOR2_X1
xU5251 n2106 n2107 n1926 VDD GND XOR2_X1
xU5252 n1916 n2091 n2107 VDD GND XOR2_X1
xU5253 n2108 n2109 n2091 VDD GND XOR2_X1
xU5254 n189 n2088 n2106 VDD GND XOR2_X1
xU5255 n2110 n2093 n2105 VDD GND XOR2_X1
xU5256 n2111 n2112 n2093 VDD GND XOR2_X1
xU5257 n2088 n2096 n2110 VDD GND XOR2_X1
xU5258 n1672 n189 n2096 VDD GND XOR2_X1
xU5259 Dout_E_3 n193 n2113 VDD GND XOR2_X1
xU5260 Dout_E_5 n2104 n1820 VDD GND XOR2_X1
xU5261 n191 n190 n2104 VDD GND XOR2_X1
xU5262 n1916 n1879 n1672 VDD GND XOR2_X1
xU5263 Dout_E_4 n2115 n2114 VDD GND XOR2_X1
xU5264 n2098 n2116 n2080 VDD GND XOR2_X1
xU5265 n186 n1763 n2116 VDD GND XOR2_X1
xU5266 n2112 n2118 n2117 VDD GND XOR2_X1
xU5267 Dout_E_1 n2120 n2119 VDD GND XOR2_X1
xU5268 n1877 n2120 n1881 VDD GND XOR2_X1
xU5269 n2108 n2121 n2098 VDD GND XOR2_X1
xU5270 n188 n1763 n2122 VDD GND XOR2_X1
xU5271 n2123 n2124 n1763 VDD GND XOR2_X1
xU5272 n1877 Dout_E_0 n1884 VDD GND XOR2_X1
xU5273 Dout_E_5 n2124 n1877 VDD GND XOR2_X1
xU5274 n2125 n2126 n1927 VDD GND XOR2_X1
xU5275 n2123 n2090 n2126 VDD GND XOR2_X1
xU5276 n2111 n2118 n2090 VDD GND XOR2_X1
xU5277 Dout_E_1 n2127 n1910 VDD GND XOR2_X1
xU5278 n1916 n2115 n1924 VDD GND XOR2_X1
xU5279 Dout_E_1 n2124 n2115 VDD GND XOR2_X1
xU5280 Dout_E_7 n1879 n2124 VDD GND XOR2_X1
xU5281 Dout_E_2 Dout_E_3 n1879 VDD GND XOR2_X1
xU5282 Dout_E_5 n193 n1916 VDD GND XOR2_X1
xU5283 n194 Dout_E_6 n2123 VDD GND XOR2_X1
xU5284 n197 n2086 n2125 VDD GND XOR2_X1
xU5285 n2121 n2109 n2086 VDD GND XOR2_X1
xU5286 Dout_E_2 n2131 n2130 VDD GND XOR2_X1
xU5287 Dout_E_3 n2131 n1911 VDD GND XOR2_X1
xU5288 n194 n197 n2131 VDD GND XOR2_X1
xU5289 n2133 n2127 n2075 VDD GND XOR2_X1
xU5290 n188 n194 n2127 VDD GND XOR2_X1
xU5291 n191 n195 n2133 VDD GND XOR2_X1
xU5292 Dout_E_3 n2120 n2132 VDD GND XOR2_X1
xU5293 n188 n196 n2120 VDD GND XOR2_X1
xU5294 n1283 n1151 n1362 VDD GND XOR2_X1
xU5295 n2134 n1348 n1151 VDD GND XOR2_X1
xU5296 n1778 n1710 n1348 VDD GND XOR2_X1
xU5297 n1216 n1831 n2134 VDD GND XOR2_X1
xU5298 n1715 n2137 n1786 VDD GND XOR2_X1
xU5299 n1153 n1797 n1283 VDD GND XOR2_X1
xU5300 n1103 n1829 n1797 VDD GND XOR2_X1
xU5301 n1648 n1719 n1829 VDD GND XOR2_X1
xU5302 n1646 n1709 n1103 VDD GND XOR2_X1
xU5303 n2143 n2144 n2137 VDD GND XOR2_X1
xU5304 n1780 n1837 n2135 VDD GND XOR2_X1
xU5305 n2146 n2144 n1837 VDD GND XOR2_X1
xU5306 n1647 n1718 n1153 VDD GND XOR2_X1
xU5307 n2152 n2153 n2147 VDD GND XOR2_X1
xU5308 n2154 n2155 n2153 VDD GND XOR2_X1
xU5309 n1783 n1835 n1832 VDD GND XOR2_X1
xU5310 n2146 n2143 n1835 VDD GND XOR2_X1
xU5311 n2160 n2161 n2152 VDD GND XOR2_X1
xU5312 n2162 n1784 n2161 VDD GND XOR2_X1
xU5313 n2163 n2164 n2157 VDD GND XOR2_X1
xU5314 n2154 n2165 n2164 VDD GND XOR2_X1
xU5315 n2167 n2168 n2159 VDD GND XOR2_X1
xU5316 n1833 n2169 n2168 VDD GND XOR2_X1
xU5317 n2170 n2171 n2166 VDD GND XOR2_X1
xU5318 n540 n2169 n2171 VDD GND XOR2_X1
xU5319 n2172 n2173 n2169 VDD GND XOR2_X1
xU5320 n2167 n2174 n2163 VDD GND XOR2_X1
xU5321 n2136 n2170 n2174 VDD GND XOR2_X1
xU5322 n2175 n2176 n2170 VDD GND XOR2_X1
xU5323 n2177 n2178 n2167 VDD GND XOR2_X1
xU5324 n2151 n2179 n2158 VDD GND XOR2_X1
xU5325 n2165 n2155 n2179 VDD GND XOR2_X1
xU5326 n2182 n2183 n2181 VDD GND XOR2_X1
xU5327 n2160 n540 n2183 VDD GND XOR2_X1
xU5328 n1833 n2136 n2138 VDD GND XOR2_X1
xU5329 n2177 n2184 n2160 VDD GND XOR2_X1
xU5330 Dout_E_80 n1784 n2185 VDD GND XOR2_X1
xU5331 n1836 Dout_E_80 n2156 VDD GND XOR2_X1
xU5332 n2182 n2186 n2180 VDD GND XOR2_X1
xU5333 n1781 n2162 n2186 VDD GND XOR2_X1
xU5334 n2176 n2187 n2162 VDD GND XOR2_X1
xU5335 Dout_E_81 n2189 n2188 VDD GND XOR2_X1
xU5336 n1836 n2189 n2141 VDD GND XOR2_X1
xU5337 Dout_E_85 n2190 n1836 VDD GND XOR2_X1
xU5338 Dout_E_85 Dout_E_87 n1781 VDD GND XOR2_X1
xU5339 n2191 n2173 n2182 VDD GND XOR2_X1
xU5340 Dout_E_83 n2193 n2192 VDD GND XOR2_X1
xU5341 n537 n2195 n2148 VDD GND XOR2_X1
xU5342 n2136 n2197 n2196 VDD GND XOR2_X1
xU5343 n2195 n2198 n2194 VDD GND XOR2_X1
xU5344 n1784 n536 n2198 VDD GND XOR2_X1
xU5345 n2193 n2190 n1784 VDD GND XOR2_X1
xU5346 n2172 n2191 n2195 VDD GND XOR2_X1
xU5347 n2200 n2201 n2199 VDD GND XOR2_X1
xU5348 Dout_E_87 Dout_E_86 n2201 VDD GND XOR2_X1
xU5349 Dout_E_86 n1830 n2149 VDD GND XOR2_X1
xU5350 Dout_E_85 n2200 n1830 VDD GND XOR2_X1
xU5351 n541 n539 n2200 VDD GND XOR2_X1
xU5352 Dout_E_84 n2203 n2202 VDD GND XOR2_X1
xU5353 n2204 n2205 n2151 VDD GND XOR2_X1
xU5354 n536 n2197 n2205 VDD GND XOR2_X1
xU5355 n2184 n2178 n2197 VDD GND XOR2_X1
xU5356 Dout_E_82 n2207 n2206 VDD GND XOR2_X1
xU5357 Dout_E_83 n2207 n2145 VDD GND XOR2_X1
xU5358 n543 n546 n2207 VDD GND XOR2_X1
xU5359 n2209 n2210 n1787 VDD GND XOR2_X1
xU5360 n541 n544 n2209 VDD GND XOR2_X1
xU5361 Dout_E_83 n2189 n2208 VDD GND XOR2_X1
xU5362 n538 n545 n2189 VDD GND XOR2_X1
xU5363 n2175 n2187 n2211 VDD GND XOR2_X1
xU5364 Dout_E_81 n2210 n2142 VDD GND XOR2_X1
xU5365 n538 n543 n2210 VDD GND XOR2_X1
xU5366 n1833 n2203 n1838 VDD GND XOR2_X1
xU5367 Dout_E_81 n2190 n2203 VDD GND XOR2_X1
xU5368 Dout_E_87 n2136 n2190 VDD GND XOR2_X1
xU5369 Dout_E_82 Dout_E_83 n2136 VDD GND XOR2_X1
xU5370 Dout_E_85 n2193 n1833 VDD GND XOR2_X1
xU5371 Dout_E_87 n2193 n2204 VDD GND XOR2_X1
xU5372 Dout_E_84 Dout_E_86 n2193 VDD GND XOR2_X1
xU5373 n777 Din_96 n2216 VDD GND XOR2_X1
xU5374 n2229 n2230 n2225 VDD GND XOR2_X1
xU5375 n2231 n2232 n2230 VDD GND XOR2_X1
xU5376 n559 n2233 n2232 VDD GND XOR2_X1
xU5377 n2234 n2235 n2229 VDD GND XOR2_X1
xU5378 n2236 n2237 n2235 VDD GND XOR2_X1
xU5379 n776 Din_95 n2240 VDD GND XOR2_X1
xU5380 n2253 n559 n2248 VDD GND XOR2_X1
xU5381 n2254 n2255 n2249 VDD GND XOR2_X1
xU5382 n2256 n2257 n2255 VDD GND XOR2_X1
xU5383 n2258 n2234 n2257 VDD GND XOR2_X1
xU5384 n2259 n2260 n2234 VDD GND XOR2_X1
xU5385 n2261 n2262 n2254 VDD GND XOR2_X1
xU5386 n775 Din_94 n2265 VDD GND XOR2_X1
xU5387 n2277 n2278 n2273 VDD GND XOR2_X1
xU5388 n2279 n2280 n2278 VDD GND XOR2_X1
xU5389 n2281 n2282 n2280 VDD GND XOR2_X1
xU5390 n2283 n2284 n2277 VDD GND XOR2_X1
xU5391 n2285 n2286 n2284 VDD GND XOR2_X1
xU5392 n774 Din_93 n2289 VDD GND XOR2_X1
xU5393 n2286 n558 n2297 VDD GND XOR2_X1
xU5394 n2302 n2303 n2298 VDD GND XOR2_X1
xU5395 n2304 n2305 n2303 VDD GND XOR2_X1
xU5396 n2306 n2307 n2305 VDD GND XOR2_X1
xU5397 n2308 n2281 n2304 VDD GND XOR2_X1
xU5398 n2309 n2310 n2302 VDD GND XOR2_X1
xU5399 n2311 n2312 n2310 VDD GND XOR2_X1
xU5400 n2313 n2314 n2309 VDD GND XOR2_X1
xU5401 n773 Din_92 n2317 VDD GND XOR2_X1
xU5402 n2330 n2331 n2326 VDD GND XOR2_X1
xU5403 n2332 n2333 n2331 VDD GND XOR2_X1
xU5404 n2334 n2335 n2333 VDD GND XOR2_X1
xU5405 n203 n2336 n2332 VDD GND XOR2_X1
xU5406 n2337 n2338 n2330 VDD GND XOR2_X1
xU5407 n2339 n2253 n2338 VDD GND XOR2_X1
xU5408 n2340 n2341 n2337 VDD GND XOR2_X1
xU5409 n772 Din_91 n2344 VDD GND XOR2_X1
xU5410 n2357 n2358 n2352 VDD GND XOR2_X1
xU5411 n2253 n2359 n2358 VDD GND XOR2_X1
xU5412 n2360 n2361 n2353 VDD GND XOR2_X1
xU5413 n2362 n2363 n2361 VDD GND XOR2_X1
xU5414 n2364 n2365 n2363 VDD GND XOR2_X1
xU5415 n2366 n2367 n2360 VDD GND XOR2_X1
xU5416 n2237 n2368 n2367 VDD GND XOR2_X1
xU5417 n2341 n2369 n2237 VDD GND XOR2_X1
xU5418 n771 Din_90 n2372 VDD GND XOR2_X1
xU5419 n2385 n2386 n2380 VDD GND XOR2_X1
xU5420 n2387 n2388 n2386 VDD GND XOR2_X1
xU5421 n2334 n2389 n2388 VDD GND XOR2_X1
xU5422 n2390 n2391 n2334 VDD GND XOR2_X1
xU5423 n2392 n2312 n2387 VDD GND XOR2_X1
xU5424 n2393 n2394 n2312 VDD GND XOR2_X1
xU5425 n2395 n2396 n2385 VDD GND XOR2_X1
xU5426 n2397 n2398 n2396 VDD GND XOR2_X1
xU5427 n2399 n2400 n2395 VDD GND XOR2_X1
xU5428 n770 Din_89 n2403 VDD GND XOR2_X1
xU5429 n2416 n2417 n2411 VDD GND XOR2_X1
xU5430 n2418 n2419 n2412 VDD GND XOR2_X1
xU5431 n2420 n2421 n2419 VDD GND XOR2_X1
xU5432 n578 n2422 n2421 VDD GND XOR2_X1
xU5433 n2423 n2424 n2418 VDD GND XOR2_X1
xU5434 n2308 n2425 n2424 VDD GND XOR2_X1
xU5435 n2426 n2394 n2423 VDD GND XOR2_X1
xU5436 n769 Din_88 n2429 VDD GND XOR2_X1
xU5437 n2442 n2369 n2437 VDD GND XOR2_X1
xU5438 n2443 n2444 n2438 VDD GND XOR2_X1
xU5439 n2445 n2446 n2444 VDD GND XOR2_X1
xU5440 n2368 n2224 n2446 VDD GND XOR2_X1
xU5441 n2447 n552 n2224 VDD GND XOR2_X1
xU5442 n2448 n2236 n2443 VDD GND XOR2_X1
xU5443 n2449 n584 n2236 VDD GND XOR2_X1
xU5444 n2450 n429 n2448 VDD GND XOR2_X1
xU5445 n768 Din_87 n2453 VDD GND XOR2_X1
xU5446 n2339 n429 n2461 VDD GND XOR2_X1
xU5447 n2466 n2467 n2462 VDD GND XOR2_X1
xU5448 n2468 n424 n2467 VDD GND XOR2_X1
xU5449 n2469 n2445 n2466 VDD GND XOR2_X1
xU5450 n239 n2470 n2445 VDD GND XOR2_X1
xU5451 n2471 n586 n2469 VDD GND XOR2_X1
xU5452 n767 Din_86 n2474 VDD GND XOR2_X1
xU5453 n2487 n2488 n2483 VDD GND XOR2_X1
xU5454 n2279 n2489 n2488 VDD GND XOR2_X1
xU5455 n549 n2490 n2489 VDD GND XOR2_X1
xU5456 n2491 n2492 n2279 VDD GND XOR2_X1
xU5457 n2493 n2494 n2487 VDD GND XOR2_X1
xU5458 n203 n2495 n2493 VDD GND XOR2_X1
xU5459 n766 Din_85 n2498 VDD GND XOR2_X1
xU5460 n2511 n2512 n2506 VDD GND XOR2_X1
xU5461 n2513 n2514 n2512 VDD GND XOR2_X1
xU5462 n577 n2515 n2514 VDD GND XOR2_X1
xU5463 n2286 n2516 n2513 VDD GND XOR2_X1
xU5464 n2517 n2518 n2511 VDD GND XOR2_X1
xU5465 n2519 n2520 n2518 VDD GND XOR2_X1
xU5466 n765 Din_84 n2523 VDD GND XOR2_X1
xU5467 n2535 n2536 n2531 VDD GND XOR2_X1
xU5468 n2537 n2538 n2536 VDD GND XOR2_X1
xU5469 n2368 n2335 n2538 VDD GND XOR2_X1
xU5470 n2366 n580 n2335 VDD GND XOR2_X1
xU5471 n2539 n2540 n2537 VDD GND XOR2_X1
xU5472 n2541 n2542 n2535 VDD GND XOR2_X1
xU5473 n2325 n2543 n2542 VDD GND XOR2_X1
xU5474 n764 Din_83 n2546 VDD GND XOR2_X1
xU5475 n2559 n2560 n2554 VDD GND XOR2_X1
xU5476 n2339 n2369 n2559 VDD GND XOR2_X1
xU5477 n2561 n2562 n2555 VDD GND XOR2_X1
xU5478 n2563 n2564 n2562 VDD GND XOR2_X1
xU5479 n2565 n2566 n2564 VDD GND XOR2_X1
xU5480 n2567 n2568 n2561 VDD GND XOR2_X1
xU5481 n2569 n2449 n2568 VDD GND XOR2_X1
xU5482 n763 Din_82 n2572 VDD GND XOR2_X1
xU5483 n2585 n2586 n2581 VDD GND XOR2_X1
xU5484 n2587 n2588 n2586 VDD GND XOR2_X1
xU5485 n2399 n2589 n2588 VDD GND XOR2_X1
xU5486 n550 n2491 n2587 VDD GND XOR2_X1
xU5487 n2543 n2590 n2585 VDD GND XOR2_X1
xU5488 n2420 n2517 n2590 VDD GND XOR2_X1
xU5489 n240 n2422 n2517 VDD GND XOR2_X1
xU5490 n427 n2391 n2422 VDD GND XOR2_X1
xU5491 n2592 n2593 n2420 VDD GND XOR2_X1
xU5492 n2594 n2595 n2593 VDD GND XOR2_X1
xU5493 n2281 n2259 n2592 VDD GND XOR2_X1
xU5494 n2596 n2597 n2543 VDD GND XOR2_X1
xU5495 n762 Din_81 n2600 VDD GND XOR2_X1
xU5496 n2613 n2614 n2609 VDD GND XOR2_X1
xU5497 n2442 n2615 n2614 VDD GND XOR2_X1
xU5498 n2616 n2417 n2615 VDD GND XOR2_X1
xU5499 n2617 n2618 n2613 VDD GND XOR2_X1
xU5500 n2520 n2591 n2617 VDD GND XOR2_X1
xU5501 n2369 n2619 n2591 VDD GND XOR2_X1
xU5502 n2416 n2490 n2520 VDD GND XOR2_X1
xU5503 n761 Din_80 n2622 VDD GND XOR2_X1
xU5504 n2635 n2636 n2630 VDD GND XOR2_X1
xU5505 n2637 n2638 n2636 VDD GND XOR2_X1
xU5506 n2639 n2425 n2638 VDD GND XOR2_X1
xU5507 n2306 n2640 n2425 VDD GND XOR2_X1
xU5508 n227 n2641 n2635 VDD GND XOR2_X1
xU5509 n2442 n2642 n2641 VDD GND XOR2_X1
xU5510 n760 Din_79 n2645 VDD GND XOR2_X1
xU5511 n2471 n2658 n2653 VDD GND XOR2_X1
xU5512 n2659 n2660 n2654 VDD GND XOR2_X1
xU5513 n2569 n2661 n2660 VDD GND XOR2_X1
xU5514 n583 n2233 n2661 VDD GND XOR2_X1
xU5515 n2662 n2468 n2659 VDD GND XOR2_X1
xU5516 n2663 n2664 n2468 VDD GND XOR2_X1
xU5517 n2665 n2666 n2664 VDD GND XOR2_X1
xU5518 n759 Din_78 n2669 VDD GND XOR2_X1
xU5519 n2682 n2666 n2677 VDD GND XOR2_X1
xU5520 n2683 n2684 n2678 VDD GND XOR2_X1
xU5521 n2685 n2686 n2684 VDD GND XOR2_X1
xU5522 n231 n2687 n2686 VDD GND XOR2_X1
xU5523 n2258 n2688 n2685 VDD GND XOR2_X1
xU5524 n2306 n2689 n2258 VDD GND XOR2_X1
xU5525 n2482 n2690 n2683 VDD GND XOR2_X1
xU5526 n2691 n2692 n2690 VDD GND XOR2_X1
xU5527 n758 Din_77 n2695 VDD GND XOR2_X1
xU5528 n2707 n2708 n2703 VDD GND XOR2_X1
xU5529 n2709 n2710 n2708 VDD GND XOR2_X1
xU5530 n420 n2711 n2710 VDD GND XOR2_X1
xU5531 n2308 n2494 n2510 VDD GND XOR2_X1
xU5532 n2712 n2713 n2707 VDD GND XOR2_X1
xU5533 n2286 n2714 n2713 VDD GND XOR2_X1
xU5534 n2715 n2716 n2286 VDD GND XOR2_X1
xU5535 n2340 n2717 n2716 VDD GND XOR2_X1
xU5536 n2718 n2719 n2715 VDD GND XOR2_X1
xU5537 n2720 n2721 n2718 VDD GND XOR2_X1
xU5538 n2722 n2723 n2712 VDD GND XOR2_X1
xU5539 n757 Din_76 n2726 VDD GND XOR2_X1
xU5540 n2565 n2739 n2734 VDD GND XOR2_X1
xU5541 n2740 n2741 n2739 VDD GND XOR2_X1
xU5542 n2742 n2743 n2741 VDD GND XOR2_X1
xU5543 n2325 n2400 n2743 VDD GND XOR2_X1
xU5544 n421 n579 n2742 VDD GND XOR2_X1
xU5545 n2744 n2745 n2740 VDD GND XOR2_X1
xU5546 n2746 n2747 n2745 VDD GND XOR2_X1
xU5547 n582 n2748 n2744 VDD GND XOR2_X1
xU5548 n2471 n2539 n2565 VDD GND XOR2_X1
xU5549 n756 Din_75 n2751 VDD GND XOR2_X1
xU5550 n2471 n2764 n2759 VDD GND XOR2_X1
xU5551 n2765 n2766 n2760 VDD GND XOR2_X1
xU5552 n2563 n2767 n2766 VDD GND XOR2_X1
xU5553 n2400 n2233 n2767 VDD GND XOR2_X1
xU5554 n2682 n2339 n2233 VDD GND XOR2_X1
xU5555 n2663 n2359 n2563 VDD GND XOR2_X1
xU5556 n2768 n2769 n2359 VDD GND XOR2_X1
xU5557 n2770 n2771 n2765 VDD GND XOR2_X1
xU5558 n2560 n2642 n2771 VDD GND XOR2_X1
xU5559 n2772 n2394 n2642 VDD GND XOR2_X1
xU5560 n755 Din_74 n2775 VDD GND XOR2_X1
xU5561 n2682 n2400 n2783 VDD GND XOR2_X1
xU5562 n2788 n2789 n2784 VDD GND XOR2_X1
xU5563 n2365 n2790 n2789 VDD GND XOR2_X1
xU5564 n2490 n2748 n2790 VDD GND XOR2_X1
xU5565 n550 n2723 n2365 VDD GND XOR2_X1
xU5566 n2306 n2336 n2384 VDD GND XOR2_X1
xU5567 n2791 n2792 n2336 VDD GND XOR2_X1
xU5568 n2340 n2768 n2306 VDD GND XOR2_X1
xU5569 n2618 n2793 n2788 VDD GND XOR2_X1
xU5570 n2794 n2580 n2793 VDD GND XOR2_X1
xU5571 n2795 n2796 n2618 VDD GND XOR2_X1
xU5572 n2797 n2711 n2796 VDD GND XOR2_X1
xU5573 n237 n2597 n2711 VDD GND XOR2_X1
xU5574 n2798 n2799 n2795 VDD GND XOR2_X1
xU5575 n754 Din_73 n2802 VDD GND XOR2_X1
xU5576 n2814 n2815 n2810 VDD GND XOR2_X1
xU5577 n419 n2816 n2815 VDD GND XOR2_X1
xU5578 n2308 n2817 n2608 VDD GND XOR2_X1
xU5579 n2449 n2417 n2814 VDD GND XOR2_X1
xU5580 n2325 n2818 n2417 VDD GND XOR2_X1
xU5581 n2540 n2723 n2449 VDD GND XOR2_X1
xU5582 n2819 n2619 n2723 VDD GND XOR2_X1
xU5583 n753 Din_72 n2822 VDD GND XOR2_X1
xU5584 n2450 n2772 n2830 VDD GND XOR2_X1
xU5585 n2835 n2836 n2831 VDD GND XOR2_X1
xU5586 n2837 n2838 n2836 VDD GND XOR2_X1
xU5587 n2839 n209 n2838 VDD GND XOR2_X1
xU5588 n2540 n2840 n2634 VDD GND XOR2_X1
xU5589 n2619 n2682 n2840 VDD GND XOR2_X1
xU5590 n2663 n2841 n2835 VDD GND XOR2_X1
xU5591 n586 n2442 n2841 VDD GND XOR2_X1
xU5592 n2519 n2341 n2442 VDD GND XOR2_X1
xU5593 n752 Din_71 n2844 VDD GND XOR2_X1
xU5594 n2747 n586 n2261 VDD GND XOR2_X1
xU5595 n2857 n2858 n2852 VDD GND XOR2_X1
xU5596 n2256 n2859 n2858 VDD GND XOR2_X1
xU5597 n2689 n2231 n2859 VDD GND XOR2_X1
xU5598 n2860 n2861 n2689 VDD GND XOR2_X1
xU5599 n2368 n2658 n2256 VDD GND XOR2_X1
xU5600 n2662 n2837 n2857 VDD GND XOR2_X1
xU5601 n2862 n2768 n2837 VDD GND XOR2_X1
xU5602 n2863 n2719 n2768 VDD GND XOR2_X1
xU5603 n2864 n2865 n2719 VDD GND XOR2_X1
xU5604 n2866 n2492 n2662 VDD GND XOR2_X1
xU5605 n751 Din_70 n2869 VDD GND XOR2_X1
xU5606 n2450 n2492 n2877 VDD GND XOR2_X1
xU5607 n2882 n2722 n2492 VDD GND XOR2_X1
xU5608 n2883 n2884 n2722 VDD GND XOR2_X1
xU5609 n2885 n2886 n2878 VDD GND XOR2_X1
xU5610 n8251 n2887 n2886 VDD GND XOR2_X1
xU5611 n2863 n2282 n2887 VDD GND XOR2_X1
xU5612 n2392 n2666 n2282 VDD GND XOR2_X1
xU5613 n2888 n2516 n2666 VDD GND XOR2_X1
xU5614 n2889 n2890 n2516 VDD GND XOR2_X1
xU5615 n2891 n424 n2885 VDD GND XOR2_X1
xU5616 n2519 n2262 n2482 VDD GND XOR2_X1
xU5617 n2892 n2307 n2262 VDD GND XOR2_X1
xU5618 n2893 n2894 n2307 VDD GND XOR2_X1
xU5619 n2325 n577 n2891 VDD GND XOR2_X1
xU5620 n2769 n2895 n2325 VDD GND XOR2_X1
xU5621 n2640 n2792 n2769 VDD GND XOR2_X1
xU5622 n750 Din_69 n2898 VDD GND XOR2_X1
xU5623 n2910 n2911 n2313 VDD GND XOR2_X1
xU5624 n2912 n2714 n2911 VDD GND XOR2_X1
xU5625 n2687 n2913 n2714 VDD GND XOR2_X1
xU5626 n2914 n2915 n2913 VDD GND XOR2_X1
xU5627 n2916 n2917 n2687 VDD GND XOR2_X1
xU5628 n2919 n593 n2918 VDD GND XOR2_X1
xU5629 n2920 n2921 n2910 VDD GND XOR2_X1
xU5630 n2922 n2923 n2920 VDD GND XOR2_X1
xU5631 n2924 n2925 n2906 VDD GND XOR2_X1
xU5632 n2926 n2927 n2925 VDD GND XOR2_X1
xU5633 n2494 n2928 n2927 VDD GND XOR2_X1
xU5634 n2929 n2930 n2494 VDD GND XOR2_X1
xU5635 n2314 n2366 n2930 VDD GND XOR2_X1
xU5636 n2931 n2285 n2314 VDD GND XOR2_X1
xU5637 n2932 n2933 n2285 VDD GND XOR2_X1
xU5638 n2936 n434 n2934 VDD GND XOR2_X1
xU5639 n2937 n2938 n2929 VDD GND XOR2_X1
xU5640 n2939 n2940 n2937 VDD GND XOR2_X1
xU5641 n2941 n2942 n2926 VDD GND XOR2_X1
xU5642 n2943 n2944 n2924 VDD GND XOR2_X1
xU5643 n2717 n2311 n2944 VDD GND XOR2_X1
xU5644 n2945 n2946 n2311 VDD GND XOR2_X1
xU5645 n2539 n2515 n2946 VDD GND XOR2_X1
xU5646 n2495 n2947 n2515 VDD GND XOR2_X1
xU5647 n2948 n2949 n2495 VDD GND XOR2_X1
xU5648 n2950 n2951 n2949 VDD GND XOR2_X1
xU5649 n245 n2954 n2952 VDD GND XOR2_X1
xU5650 n2955 n2956 n2945 VDD GND XOR2_X1
xU5651 n2957 n2958 n2955 VDD GND XOR2_X1
xU5652 n2959 n8251 n2717 VDD GND XOR2_X1
xU5654 n2965 n563 n2963 VDD GND XOR2_X1
xU5655 n2819 n2861 n2943 VDD GND XOR2_X1
xU5656 n2966 n2967 n2861 VDD GND XOR2_X1
xU5657 n749 Din_68 n2970 VDD GND XOR2_X1
xU5658 n2691 n2942 n2978 VDD GND XOR2_X1
xU5659 n2983 n2984 n2979 VDD GND XOR2_X1
xU5660 n2985 n2986 n2984 VDD GND XOR2_X1
xU5661 n2663 n2770 n2986 VDD GND XOR2_X1
xU5662 n2912 n2791 n2770 VDD GND XOR2_X1
xU5663 n2253 n2747 n2663 VDD GND XOR2_X1
xU5664 n2987 n2988 n2983 VDD GND XOR2_X1
xU5665 n2895 n2738 n2988 VDD GND XOR2_X1
xU5666 n2283 n2640 n2987 VDD GND XOR2_X1
xU5667 n748 Din_67 n2991 VDD GND XOR2_X1
xU5668 n2819 n2362 n2999 VDD GND XOR2_X1
xU5669 n2567 n2637 n2362 VDD GND XOR2_X1
xU5670 n2569 n2747 n2637 VDD GND XOR2_X1
xU5671 n3004 n3005 n2747 VDD GND XOR2_X1
xU5672 n3006 n2916 n3005 VDD GND XOR2_X1
xU5673 n593 n3009 n3007 VDD GND XOR2_X1
xU5674 n2691 n2748 n2567 VDD GND XOR2_X1
xU5675 n3012 n3013 n3000 VDD GND XOR2_X1
xU5676 n2985 n3014 n3013 VDD GND XOR2_X1
xU5677 n2839 n2764 n3014 VDD GND XOR2_X1
xU5678 n2619 n2364 n2764 VDD GND XOR2_X1
xU5679 n3015 n3016 n2364 VDD GND XOR2_X1
xU5680 n2596 n2470 n3016 VDD GND XOR2_X1
xU5681 n2394 n556 n2839 VDD GND XOR2_X1
xU5682 n2860 n2959 n2640 VDD GND XOR2_X1
xU5683 n2447 n2369 n2394 VDD GND XOR2_X1
xU5684 n2340 n2399 n2985 VDD GND XOR2_X1
xU5685 n559 n2862 n2340 VDD GND XOR2_X1
xU5686 n2560 n3025 n3012 VDD GND XOR2_X1
xU5687 n2231 n2368 n3025 VDD GND XOR2_X1
xU5688 n2339 n2471 n2368 VDD GND XOR2_X1
xU5689 n3026 n3027 n2471 VDD GND XOR2_X1
xU5690 n3028 n2950 n3027 VDD GND XOR2_X1
xU5691 n245 n3031 n3029 VDD GND XOR2_X1
xU5692 n2932 n3034 n2339 VDD GND XOR2_X1
xU5693 n2595 n3035 n3034 VDD GND XOR2_X1
xU5694 n434 n3040 n3038 VDD GND XOR2_X1
xU5695 n2450 n2253 n2231 VDD GND XOR2_X1
xU5696 n2961 n3041 n2253 VDD GND XOR2_X1
xU5697 n3042 n3043 n3041 VDD GND XOR2_X1
xU5698 n567 n3048 n3046 VDD GND XOR2_X1
xU5699 n3049 n3050 n2560 VDD GND XOR2_X1
xU5700 n2390 n2260 n3050 VDD GND XOR2_X1
xU5701 n747 Din_66 n3053 VDD GND XOR2_X1
xU5702 n2450 n2399 n3061 VDD GND XOR2_X1
xU5703 n2748 n2941 n2399 VDD GND XOR2_X1
xU5704 n3068 n3069 n3062 VDD GND XOR2_X1
xU5705 n2816 n3070 n3069 VDD GND XOR2_X1
xU5706 n2818 n2566 n3070 VDD GND XOR2_X1
xU5707 n2580 n2357 n2566 VDD GND XOR2_X1
xU5708 n2447 n2791 n2357 VDD GND XOR2_X1
xU5709 n2519 n2541 n2580 VDD GND XOR2_X1
xU5710 n2390 n3074 n2541 VDD GND XOR2_X1
xU5711 n2366 n2260 n2519 VDD GND XOR2_X1
xU5712 n2281 n2938 n2260 VDD GND XOR2_X1
xU5713 n2594 n3078 n2938 VDD GND XOR2_X1
xU5714 Dout_E_49 n3082 n3080 VDD GND XOR2_X1
xU5715 n429 n2259 n2366 VDD GND XOR2_X1
xU5716 n3042 n3085 n2818 VDD GND XOR2_X1
xU5717 n2665 n2865 n3085 VDD GND XOR2_X1
xU5718 n3086 n3087 n3019 VDD GND XOR2_X1
xU5719 n3089 n564 n2965 VDD GND XOR2_X1
xU5720 n3090 n3091 n2816 VDD GND XOR2_X1
xU5721 n3092 n2709 n3091 VDD GND XOR2_X1
xU5722 n2392 n2688 n2709 VDD GND XOR2_X1
xU5723 n2682 n558 n2392 VDD GND XOR2_X1
xU5724 n2539 n2470 n2682 VDD GND XOR2_X1
xU5725 n2490 n2956 n2470 VDD GND XOR2_X1
xU5726 n2798 n3093 n2956 VDD GND XOR2_X1
xU5727 Dout_E_9 n3097 n3095 VDD GND XOR2_X1
xU5728 n2658 n239 n2539 VDD GND XOR2_X1
xU5729 n3100 n2941 n3090 VDD GND XOR2_X1
xU5730 n3101 n2639 n3100 VDD GND XOR2_X1
xU5731 n2400 n3102 n3068 VDD GND XOR2_X1
xU5732 n2819 n2895 n3102 VDD GND XOR2_X1
xU5733 n2596 n237 n2400 VDD GND XOR2_X1
xU5734 n746 Din_65 n3108 VDD GND XOR2_X1
xU5735 n2691 n2794 n2616 VDD GND XOR2_X1
xU5736 n3120 n3092 n2794 VDD GND XOR2_X1
xU5737 n2692 n3004 n3092 VDD GND XOR2_X1
xU5738 n579 n2915 n2692 VDD GND XOR2_X1
xU5739 n2883 n2922 n2942 VDD GND XOR2_X1
xU5740 n2856 n3128 n3120 VDD GND XOR2_X1
xU5741 n2746 n2941 n2691 VDD GND XOR2_X1
xU5742 n2884 n2923 n2941 VDD GND XOR2_X1
xU5743 n3130 n3131 n3116 VDD GND XOR2_X1
xU5744 n2928 n3132 n3131 VDD GND XOR2_X1
xU5745 n2817 n2772 n3132 VDD GND XOR2_X1
xU5746 n584 n2819 n2772 VDD GND XOR2_X1
xU5747 n2882 n2914 n2746 VDD GND XOR2_X1
xU5748 n3010 n3123 n3121 VDD GND XOR2_X1
xU5749 n2283 n2398 n2817 VDD GND XOR2_X1
xU5750 n2595 n3140 n2398 VDD GND XOR2_X1
xU5751 n2866 n3078 n3140 VDD GND XOR2_X1
xU5752 n3142 n3143 n3023 VDD GND XOR2_X1
xU5753 n3144 n3077 n3142 VDD GND XOR2_X1
xU5754 n3049 n2391 n2283 VDD GND XOR2_X1
xU5755 n2893 n2939 n2391 VDD GND XOR2_X1
xU5756 n3149 n3143 n3079 VDD GND XOR2_X1
xU5757 n3150 n3076 n3143 VDD GND XOR2_X1
xU5758 n3151 n3152 n3149 VDD GND XOR2_X1
xU5759 n2341 n427 n3049 VDD GND XOR2_X1
xU5760 n2894 n2940 n3074 VDD GND XOR2_X1
xU5761 n3152 n3150 n3081 VDD GND XOR2_X1
xU5762 n2892 n2931 n2341 VDD GND XOR2_X1
xU5763 n3144 n3150 n3141 VDD GND XOR2_X1
xU5764 n3158 n3159 n3153 VDD GND XOR2_X1
xU5765 n3160 n3161 n3159 VDD GND XOR2_X1
xU5766 n3036 n3083 n3145 VDD GND XOR2_X1
xU5767 n3165 n3166 n3158 VDD GND XOR2_X1
xU5768 n3146 n3167 n3166 VDD GND XOR2_X1
xU5769 n3169 n2389 n2928 VDD GND XOR2_X1
xU5770 n2491 n2863 n2389 VDD GND XOR2_X1
xU5771 n570 n3048 n3170 VDD GND XOR2_X1
xU5772 n2450 n2308 n2491 VDD GND XOR2_X1
xU5773 n3152 n3144 n3083 VDD GND XOR2_X1
xU5774 n3154 n3173 n3164 VDD GND XOR2_X1
xU5775 n3160 n3174 n3173 VDD GND XOR2_X1
xU5776 n3167 n3177 n3175 VDD GND XOR2_X1
xU5777 n435 n3178 n3177 VDD GND XOR2_X1
xU5778 n3179 n3180 n3167 VDD GND XOR2_X1
xU5779 n3181 n3182 n3154 VDD GND XOR2_X1
xU5780 n3040 n3183 n3182 VDD GND XOR2_X1
xU5781 n3165 n3184 n3176 VDD GND XOR2_X1
xU5782 n3185 n3178 n3184 VDD GND XOR2_X1
xU5783 n3186 n3187 n3178 VDD GND XOR2_X1
xU5784 n3188 n3189 n3165 VDD GND XOR2_X1
xU5785 n3163 n3190 n3168 VDD GND XOR2_X1
xU5786 n3174 n3161 n3190 VDD GND XOR2_X1
xU5787 n3192 n3193 n3172 VDD GND XOR2_X1
xU5788 n3146 n3194 n3192 VDD GND XOR2_X1
xU5789 n3193 n3195 n3191 VDD GND XOR2_X1
xU5790 n3040 n3196 n3195 VDD GND XOR2_X1
xU5791 n3186 n3197 n3193 VDD GND XOR2_X1
xU5792 Dout_E_52 n3199 n3198 VDD GND XOR2_X1
xU5793 n3201 n3202 n3200 VDD GND XOR2_X1
xU5794 n3037 n3181 n3202 VDD GND XOR2_X1
xU5795 n3180 n3203 n3181 VDD GND XOR2_X1
xU5796 Dout_E_49 n3205 n3204 VDD GND XOR2_X1
xU5797 n3082 n3205 n3155 VDD GND XOR2_X1
xU5798 Dout_E_53 Dout_E_55 n3037 VDD GND XOR2_X1
xU5799 n2936 n3206 n3157 VDD GND XOR2_X1
xU5800 n3183 n3201 n3206 VDD GND XOR2_X1
xU5801 n3197 n3187 n3201 VDD GND XOR2_X1
xU5802 Dout_E_51 n439 n3207 VDD GND XOR2_X1
xU5803 n3209 n3210 n3208 VDD GND XOR2_X1
xU5804 Dout_E_55 Dout_E_54 n3210 VDD GND XOR2_X1
xU5805 Dout_E_54 n3075 n3147 VDD GND XOR2_X1
xU5806 Dout_E_53 n3209 n3075 VDD GND XOR2_X1
xU5807 n436 n434 n3209 VDD GND XOR2_X1
xU5808 n3188 n3211 n3183 VDD GND XOR2_X1
xU5809 n433 n3040 n3212 VDD GND XOR2_X1
xU5810 n3213 n3214 n3040 VDD GND XOR2_X1
xU5811 n3082 Dout_E_48 n3148 VDD GND XOR2_X1
xU5812 Dout_E_53 n3214 n3082 VDD GND XOR2_X1
xU5813 n438 n3146 n2936 VDD GND XOR2_X1
xU5814 n3215 n3216 n3163 VDD GND XOR2_X1
xU5815 n3196 n3194 n3216 VDD GND XOR2_X1
xU5816 n3211 n3189 n3194 VDD GND XOR2_X1
xU5817 Dout_E_50 n3218 n3217 VDD GND XOR2_X1
xU5818 Dout_E_51 n3218 n3162 VDD GND XOR2_X1
xU5819 n440 n443 n3218 VDD GND XOR2_X1
xU5820 n3220 n3221 n3024 VDD GND XOR2_X1
xU5821 n436 n441 n3220 VDD GND XOR2_X1
xU5822 Dout_E_51 n3205 n3219 VDD GND XOR2_X1
xU5823 n433 n442 n3205 VDD GND XOR2_X1
xU5824 n3179 n3203 n3196 VDD GND XOR2_X1
xU5825 Dout_E_49 n3221 n3156 VDD GND XOR2_X1
xU5826 n433 n440 n3221 VDD GND XOR2_X1
xU5827 n438 n3199 n3084 VDD GND XOR2_X1
xU5828 Dout_E_49 n3214 n3199 VDD GND XOR2_X1
xU5829 Dout_E_55 n3146 n3214 VDD GND XOR2_X1
xU5830 Dout_E_50 Dout_E_51 n3146 VDD GND XOR2_X1
xU5831 n441 n439 n3185 VDD GND XOR2_X1
xU5832 n443 n3213 n3215 VDD GND XOR2_X1
xU5833 n440 Dout_E_54 n3213 VDD GND XOR2_X1
xU5834 n2569 n582 n2450 VDD GND XOR2_X1
xU5835 n2856 n583 n2912 VDD GND XOR2_X1
xU5836 n3225 n3226 n3123 VDD GND XOR2_X1
xU5837 n588 n3136 n3133 VDD GND XOR2_X1
xU5838 n2688 n2921 n2569 VDD GND XOR2_X1
xU5839 n3101 n3128 n2921 VDD GND XOR2_X1
xU5840 n3226 n3230 n3136 VDD GND XOR2_X1
xU5841 n3232 n3233 n3229 VDD GND XOR2_X1
xU5842 n3234 n3235 n3233 VDD GND XOR2_X1
xU5843 n3008 n581 n3126 VDD GND XOR2_X1
xU5844 n3238 n3239 n3232 VDD GND XOR2_X1
xU5845 n590 n3009 n3239 VDD GND XOR2_X1
xU5846 n3225 n3230 n3243 VDD GND XOR2_X1
xU5847 n3241 n3245 n3237 VDD GND XOR2_X1
xU5848 n3234 n3246 n3245 VDD GND XOR2_X1
xU5849 n3249 n3250 n3247 VDD GND XOR2_X1
xU5850 n3251 n3252 n3249 VDD GND XOR2_X1
xU5851 n3253 n3254 n3241 VDD GND XOR2_X1
xU5852 n3122 n3250 n3254 VDD GND XOR2_X1
xU5853 n3255 n3256 n3250 VDD GND XOR2_X1
xU5854 n3257 n3258 n3248 VDD GND XOR2_X1
xU5855 n3236 n3253 n3258 VDD GND XOR2_X1
xU5856 n3259 n3260 n3253 VDD GND XOR2_X1
xU5857 n592 n3251 n3257 VDD GND XOR2_X1
xU5858 n3228 n3261 n3240 VDD GND XOR2_X1
xU5859 n3246 n3235 n3261 VDD GND XOR2_X1
xU5860 n3252 n3263 n3244 VDD GND XOR2_X1
xU5861 n3264 n3238 n3263 VDD GND XOR2_X1
xU5862 n3259 n3265 n3238 VDD GND XOR2_X1
xU5863 n591 n3009 n3266 VDD GND XOR2_X1
xU5864 n3124 Dout_E_96 n3127 VDD GND XOR2_X1
xU5865 n2919 n592 n3252 VDD GND XOR2_X1
xU5866 n3236 n3122 n2919 VDD GND XOR2_X1
xU5867 n3268 n3269 n3262 VDD GND XOR2_X1
xU5868 n3011 n590 n3269 VDD GND XOR2_X1
xU5869 n3256 n3271 n3270 VDD GND XOR2_X1
xU5870 Dout_E_97 n3273 n3272 VDD GND XOR2_X1
xU5871 n3124 n3273 n3129 VDD GND XOR2_X1
xU5872 Dout_E_103 Dout_E_101 n3011 VDD GND XOR2_X1
xU5873 n3267 n3264 n3268 VDD GND XOR2_X1
xU5874 Dout_E_99 n596 n3274 VDD GND XOR2_X1
xU5875 Dout_E_101 n3275 n3067 VDD GND XOR2_X1
xU5876 n3277 n3278 n3231 VDD GND XOR2_X1
xU5877 n3122 n3279 n3277 VDD GND XOR2_X1
xU5878 n589 n3280 n3276 VDD GND XOR2_X1
xU5879 n3278 n3009 n3280 VDD GND XOR2_X1
xU5880 n3281 n3282 n3009 VDD GND XOR2_X1
xU5881 n3251 n3264 n3278 VDD GND XOR2_X1
xU5882 Dout_E_103 n3284 n3283 VDD GND XOR2_X1
xU5883 Dout_E_101 n3284 n3125 VDD GND XOR2_X1
xU5884 Dout_E_102 n3275 n3284 VDD GND XOR2_X1
xU5885 n594 n593 n3275 VDD GND XOR2_X1
xU5886 Dout_E_100 n3286 n3285 VDD GND XOR2_X1
xU5887 n3288 n3289 n3228 VDD GND XOR2_X1
xU5888 n3281 n3287 n3289 VDD GND XOR2_X1
xU5889 n3255 n3271 n3287 VDD GND XOR2_X1
xU5890 Dout_E_97 n3290 n3135 VDD GND XOR2_X1
xU5891 n3236 n3286 n3224 VDD GND XOR2_X1
xU5892 Dout_E_97 n3282 n3286 VDD GND XOR2_X1
xU5893 Dout_E_101 n596 n3236 VDD GND XOR2_X1
xU5894 n597 Dout_E_102 n3281 VDD GND XOR2_X1
xU5895 n600 n3279 n3288 VDD GND XOR2_X1
xU5896 n3265 n3260 n3279 VDD GND XOR2_X1
xU5897 Dout_E_99 n3294 n3137 VDD GND XOR2_X1
xU5898 Dout_E_98 n3294 n3293 VDD GND XOR2_X1
xU5899 n597 n600 n3294 VDD GND XOR2_X1
xU5900 Dout_E_99 n3273 n3295 VDD GND XOR2_X1
xU5901 n599 n591 n3273 VDD GND XOR2_X1
xU5902 n3296 n3290 n3134 VDD GND XOR2_X1
xU5903 n597 n591 n3290 VDD GND XOR2_X1
xU5904 n594 n598 n3296 VDD GND XOR2_X1
xU5905 Dout_E_97 n3124 n3242 VDD GND XOR2_X1
xU5906 Dout_E_101 n3282 n3124 VDD GND XOR2_X1
xU5907 Dout_E_103 n3122 n3282 VDD GND XOR2_X1
xU5908 Dout_E_98 Dout_E_99 n3122 VDD GND XOR2_X1
xU5909 n2447 n2416 n3169 VDD GND XOR2_X1
xU5910 n3300 n3301 n3088 VDD GND XOR2_X1
xU5911 n3087 n3073 n3300 VDD GND XOR2_X1
xU5912 n2426 n3302 n3130 VDD GND XOR2_X1
xU5913 n2393 n2397 n3302 VDD GND XOR2_X1
xU5914 n3303 n3042 n2397 VDD GND XOR2_X1
xU5915 n3044 n3297 n3021 VDD GND XOR2_X1
xU5916 n2864 n2862 n3303 VDD GND XOR2_X1
xU5917 n3304 n3087 n3297 VDD GND XOR2_X1
xU5918 n2895 n2792 n2393 VDD GND XOR2_X1
xU5919 n2967 n2720 n2792 VDD GND XOR2_X1
xU5920 n3086 n3304 n3171 VDD GND XOR2_X1
xU5921 n2966 n2721 n2895 VDD GND XOR2_X1
xU5922 n3312 n3313 n3305 VDD GND XOR2_X1
xU5923 n3314 n3315 n3313 VDD GND XOR2_X1
xU5924 n3317 n3301 n3307 VDD GND XOR2_X1
xU5925 n3086 n3072 n3301 VDD GND XOR2_X1
xU5926 n3319 n3320 n3312 VDD GND XOR2_X1
xU5927 n3321 n3322 n3320 VDD GND XOR2_X1
xU5928 n3324 n3325 n3318 VDD GND XOR2_X1
xU5929 n3314 n3326 n3325 VDD GND XOR2_X1
xU5930 n3329 n3330 n3327 VDD GND XOR2_X1
xU5931 n3331 n3332 n3330 VDD GND XOR2_X1
xU5932 n3333 n3334 n3329 VDD GND XOR2_X1
xU5933 n3308 n3304 n3317 VDD GND XOR2_X1
xU5934 n3336 n3337 n3328 VDD GND XOR2_X1
xU5935 n3338 n3339 n3324 VDD GND XOR2_X1
xU5936 n3333 n3319 n3339 VDD GND XOR2_X1
xU5937 n3340 n3334 n3319 VDD GND XOR2_X1
xU5938 n3311 n3341 n3335 VDD GND XOR2_X1
xU5939 n3315 n3326 n3341 VDD GND XOR2_X1
xU5940 n3343 n3336 n3306 VDD GND XOR2_X1
xU5941 n3344 n3345 n3336 VDD GND XOR2_X1
xU5942 n3346 n3347 n3342 VDD GND XOR2_X1
xU5943 n3322 n3332 n3347 VDD GND XOR2_X1
xU5944 n3348 n3344 n3332 VDD GND XOR2_X1
xU5945 n568 n3048 n3349 VDD GND XOR2_X1
xU5946 n3350 n3351 n3346 VDD GND XOR2_X1
xU5947 n3343 n3337 n3323 VDD GND XOR2_X1
xU5948 n3340 n3331 n3337 VDD GND XOR2_X1
xU5949 n3089 n3353 n3331 VDD GND XOR2_X1
xU5950 n3322 n3355 n3354 VDD GND XOR2_X1
xU5951 n561 n567 n3355 VDD GND XOR2_X1
xU5952 n3298 Dout_E_88 n3316 VDD GND XOR2_X1
xU5953 n3333 n3356 n3343 VDD GND XOR2_X1
xU5954 n3350 n3357 n3356 VDD GND XOR2_X1
xU5955 n3358 n3359 n3352 VDD GND XOR2_X1
xU5956 n3334 n3353 n3359 VDD GND XOR2_X1
xU5957 n566 n567 n3360 VDD GND XOR2_X1
xU5958 Dout_E_89 n3361 n3071 VDD GND XOR2_X1
xU5959 Dout_E_89 n3363 n3362 VDD GND XOR2_X1
xU5960 n3298 n3363 n3309 VDD GND XOR2_X1
xU5961 n3322 Dout_E_93 n3298 VDD GND XOR2_X1
xU5962 n3364 n3365 n3358 VDD GND XOR2_X1
xU5963 n3367 n3368 n3366 VDD GND XOR2_X1
xU5964 Dout_E_95 Dout_E_90 n3368 VDD GND XOR2_X1
xU5965 n3367 n3361 n3310 VDD GND XOR2_X1
xU5966 Dout_E_94 Dout_E_89 n3367 VDD GND XOR2_X1
xU5967 n570 Dout_E_95 n3045 VDD GND XOR2_X1
xU5968 n3369 n3338 n3311 VDD GND XOR2_X1
xU5969 n3348 n3345 n3338 VDD GND XOR2_X1
xU5970 Dout_E_90 n3371 n3370 VDD GND XOR2_X1
xU5971 Dout_E_91 n3371 n3022 VDD GND XOR2_X1
xU5972 n568 n572 n3371 VDD GND XOR2_X1
xU5973 n3048 n3089 n3374 VDD GND XOR2_X1
xU5974 n570 n567 n3089 VDD GND XOR2_X1
xU5975 n3322 n563 n3048 VDD GND XOR2_X1
xU5976 Dout_E_95 n564 n3322 VDD GND XOR2_X1
xU5977 n565 Dout_E_91 n3333 VDD GND XOR2_X1
xU5978 n572 n3321 n3369 VDD GND XOR2_X1
xU5979 n3357 n3351 n3321 VDD GND XOR2_X1
xU5980 n3365 n3375 n3351 VDD GND XOR2_X1
xU5981 Dout_E_92 Dout_E_94 n3375 VDD GND XOR2_X1
xU5982 Dout_E_89 n3376 n3020 VDD GND XOR2_X1
xU5983 n3361 n3376 n3299 VDD GND XOR2_X1
xU5984 n561 n568 n3376 VDD GND XOR2_X1
xU5985 Dout_E_90 Dout_E_93 n3361 VDD GND XOR2_X1
xU5986 Dout_E_91 n3363 n3377 VDD GND XOR2_X1
xU5987 n561 n571 n3363 VDD GND XOR2_X1
xU5988 n203 n2589 n2426 VDD GND XOR2_X1
xU5989 n3378 n2797 n2589 VDD GND XOR2_X1
xU5990 n3026 n2948 n2797 VDD GND XOR2_X1
xU5991 n2658 n3093 n3378 VDD GND XOR2_X1
xU5992 n3381 n3382 n3017 VDD GND XOR2_X1
xU5993 n3383 n3105 n3382 VDD GND XOR2_X1
xU5994 n3015 n2597 n2738 VDD GND XOR2_X1
xU5995 n2889 n2957 n2597 VDD GND XOR2_X1
xU5996 n3381 n3386 n3094 VDD GND XOR2_X1
xU5997 n3387 n3388 n3386 VDD GND XOR2_X1
xU5998 n3389 n3104 n3381 VDD GND XOR2_X1
xU5999 n2540 n237 n3015 VDD GND XOR2_X1
xU6000 n2890 n2958 n3390 VDD GND XOR2_X1
xU6001 n3387 n3389 n3096 VDD GND XOR2_X1
xU6002 n2888 n2947 n2540 VDD GND XOR2_X1
xU6003 n3383 n3389 n3380 VDD GND XOR2_X1
xU6004 n3395 n3396 n3391 VDD GND XOR2_X1
xU6005 n3032 n3098 n3379 VDD GND XOR2_X1
xU6006 n3383 n3387 n3098 VDD GND XOR2_X1
xU6007 n241 n3405 n3402 VDD GND XOR2_X1
xU6008 n3398 n3406 n3405 VDD GND XOR2_X1
xU6009 n3408 n3409 n3401 VDD GND XOR2_X1
xU6010 n3410 n3411 n3409 VDD GND XOR2_X1
xU6011 n3412 n3413 n3408 VDD GND XOR2_X1
xU6012 n3414 n3415 n3407 VDD GND XOR2_X1
xU6013 n3413 n3416 n3414 VDD GND XOR2_X1
xU6014 n3418 n3419 n3417 VDD GND XOR2_X1
xU6015 n3031 n3420 n3419 VDD GND XOR2_X1
xU6016 n242 n3421 n3396 VDD GND XOR2_X1
xU6017 n3422 n3411 n3421 VDD GND XOR2_X1
xU6018 n3423 n3424 n3411 VDD GND XOR2_X1
xU6019 n3425 n3426 n3415 VDD GND XOR2_X1
xU6020 n3404 n3427 n3400 VDD GND XOR2_X1
xU6021 n3406 n3397 n3427 VDD GND XOR2_X1
xU6022 n3429 n3430 n3403 VDD GND XOR2_X1
xU6023 n3422 n3431 n3430 VDD GND XOR2_X1
xU6024 n3432 n3433 n3428 VDD GND XOR2_X1
xU6025 n3031 n3431 n3433 VDD GND XOR2_X1
xU6026 n3413 n244 n3431 VDD GND XOR2_X1
xU6027 Dout_E_12 n3435 n3434 VDD GND XOR2_X1
xU6028 n3416 n3437 n3394 VDD GND XOR2_X1
xU6029 n3438 n3420 n3437 VDD GND XOR2_X1
xU6030 n3423 n3439 n3420 VDD GND XOR2_X1
xU6031 n243 n3031 n3440 VDD GND XOR2_X1
xU6032 n3441 n3442 n3031 VDD GND XOR2_X1
xU6033 n3097 Dout_E_8 n3385 VDD GND XOR2_X1
xU6034 n2954 n3412 n3416 VDD GND XOR2_X1
xU6035 n3410 n247 n2954 VDD GND XOR2_X1
xU6036 n3443 n3444 n3436 VDD GND XOR2_X1
xU6037 n3033 n3418 n3444 VDD GND XOR2_X1
xU6038 n3426 n3445 n3418 VDD GND XOR2_X1
xU6039 Dout_E_9 n3447 n3446 VDD GND XOR2_X1
xU6040 n3097 n3447 n3392 VDD GND XOR2_X1
xU6041 Dout_E_13 n3442 n3097 VDD GND XOR2_X1
xU6042 Dout_E_13 Dout_E_15 n3033 VDD GND XOR2_X1
xU6043 n244 n3412 n3443 VDD GND XOR2_X1
xU6044 Dout_E_11 n251 n3448 VDD GND XOR2_X1
xU6045 Dout_E_9 n3449 n3103 VDD GND XOR2_X1
xU6046 n3451 n3452 n3450 VDD GND XOR2_X1
xU6047 n3449 n3451 n3384 VDD GND XOR2_X1
xU6048 n254 n245 n3451 VDD GND XOR2_X1
xU6049 n3453 n3454 n3404 VDD GND XOR2_X1
xU6050 n3429 n3432 n3454 VDD GND XOR2_X1
xU6051 n3425 n3445 n3432 VDD GND XOR2_X1
xU6052 Dout_E_9 n3455 n3393 VDD GND XOR2_X1
xU6053 n250 n3435 n3099 VDD GND XOR2_X1
xU6054 Dout_E_9 n3442 n3435 VDD GND XOR2_X1
xU6055 n255 n3422 n3442 VDD GND XOR2_X1
xU6056 n248 Dout_E_11 n3422 VDD GND XOR2_X1
xU6057 n253 n251 n3410 VDD GND XOR2_X1
xU6058 n3439 n3424 n3429 VDD GND XOR2_X1
xU6059 Dout_E_11 n3459 n3399 VDD GND XOR2_X1
xU6060 Dout_E_15 Dout_E_12 n3459 VDD GND XOR2_X1
xU6061 Dout_E_12 n3452 n3458 VDD GND XOR2_X1
xU6062 n248 n255 n3452 VDD GND XOR2_X1
xU6063 Dout_E_11 n3447 n3460 VDD GND XOR2_X1
xU6064 n254 n243 n3447 VDD GND XOR2_X1
xU6065 n3449 n3455 n3018 VDD GND XOR2_X1
xU6066 n252 n243 n3455 VDD GND XOR2_X1
xU6067 Dout_E_10 Dout_E_13 n3449 VDD GND XOR2_X1
xU6068 n255 n3441 n3453 VDD GND XOR2_X1
xU6069 n252 Dout_E_14 n3441 VDD GND XOR2_X1
xU6070 n745 Din_64 n3463 VDD GND XOR2_X1
xU6071 n3476 n455 n3471 VDD GND XOR2_X1
xU6072 n3477 n3478 n3472 VDD GND XOR2_X1
xU6073 n3479 n3480 n3478 VDD GND XOR2_X1
xU6074 n3481 n3482 n3480 VDD GND XOR2_X1
xU6075 n3483 n3484 n3477 VDD GND XOR2_X1
xU6076 n3485 n3486 n3484 VDD GND XOR2_X1
xU6077 n744 Din_63 n3489 VDD GND XOR2_X1
xU6078 n3502 n3503 n3497 VDD GND XOR2_X1
xU6079 n3504 n3505 n3503 VDD GND XOR2_X1
xU6080 n3506 n3507 n3505 VDD GND XOR2_X1
xU6081 n3508 n3483 n3502 VDD GND XOR2_X1
xU6082 n3509 n3510 n3483 VDD GND XOR2_X1
xU6083 n297 n3511 n3508 VDD GND XOR2_X1
xU6084 n743 Din_62 n3514 VDD GND XOR2_X1
xU6085 n3526 n3527 n3522 VDD GND XOR2_X1
xU6086 n3528 n3529 n3527 VDD GND XOR2_X1
xU6087 n3530 n3531 n3529 VDD GND XOR2_X1
xU6088 n471 n3532 n3526 VDD GND XOR2_X1
xU6089 n262 n3533 n3532 VDD GND XOR2_X1
xU6090 n742 Din_61 n3536 VDD GND XOR2_X1
xU6091 n3548 n3549 n3544 VDD GND XOR2_X1
xU6092 n3550 n3551 n3549 VDD GND XOR2_X1
xU6093 n3552 n3553 n3551 VDD GND XOR2_X1
xU6094 n3531 n3554 n3550 VDD GND XOR2_X1
xU6095 n3555 n3556 n3548 VDD GND XOR2_X1
xU6096 n472 n3557 n3556 VDD GND XOR2_X1
xU6097 n3558 n3559 n3555 VDD GND XOR2_X1
xU6098 n741 Din_60 n3562 VDD GND XOR2_X1
xU6099 n3575 n3576 n3571 VDD GND XOR2_X1
xU6100 n452 n3577 n3576 VDD GND XOR2_X1
xU6101 n3578 n3579 n3577 VDD GND XOR2_X1
xU6102 n3580 n3581 n3579 VDD GND XOR2_X1
xU6103 n478 n3582 n3581 VDD GND XOR2_X1
xU6104 n3583 n3584 n3578 VDD GND XOR2_X1
xU6105 n3485 n3585 n3584 VDD GND XOR2_X1
xU6106 n3586 n298 n3575 VDD GND XOR2_X1
xU6107 n740 Din_59 n3589 VDD GND XOR2_X1
xU6108 n3602 n3603 n3597 VDD GND XOR2_X1
xU6109 n3604 n456 n3602 VDD GND XOR2_X1
xU6110 n3605 n3606 n3598 VDD GND XOR2_X1
xU6111 n3607 n3608 n3606 VDD GND XOR2_X1
xU6112 n3486 n3609 n3608 VDD GND XOR2_X1
xU6113 n3585 n3610 n3486 VDD GND XOR2_X1
xU6114 n3611 n3612 n3605 VDD GND XOR2_X1
xU6115 n3613 n3614 n3612 VDD GND XOR2_X1
xU6116 n739 Din_58 n3617 VDD GND XOR2_X1
xU6117 n3586 n3553 n3625 VDD GND XOR2_X1
xU6118 n3630 n3631 n3626 VDD GND XOR2_X1
xU6119 n3632 n3633 n3631 VDD GND XOR2_X1
xU6120 n3583 n3559 n3633 VDD GND XOR2_X1
xU6121 n3634 n3635 n3630 VDD GND XOR2_X1
xU6122 n3636 n3637 n3635 VDD GND XOR2_X1
xU6123 n738 Din_57 n3640 VDD GND XOR2_X1
xU6124 n3653 n3654 n3649 VDD GND XOR2_X1
xU6125 n601 n3655 n3654 VDD GND XOR2_X1
xU6126 n474 n3656 n3655 VDD GND XOR2_X1
xU6127 n3559 n3657 n3653 VDD GND XOR2_X1
xU6128 n3476 n3658 n3657 VDD GND XOR2_X1
xU6129 n455 n3659 n3559 VDD GND XOR2_X1
xU6130 n737 Din_56 n3662 VDD GND XOR2_X1
xU6131 n3675 n3676 n3671 VDD GND XOR2_X1
xU6132 n3476 n3677 n3676 VDD GND XOR2_X1
xU6133 n3678 n3679 n3677 VDD GND XOR2_X1
xU6134 n3680 n3681 n3675 VDD GND XOR2_X1
xU6135 n3682 n296 n3681 VDD GND XOR2_X1
xU6136 n736 Din_55 n3685 VDD GND XOR2_X1
xU6137 n297 n3698 n3693 VDD GND XOR2_X1
xU6138 n3699 n3700 n3694 VDD GND XOR2_X1
xU6139 n3701 n3702 n3700 VDD GND XOR2_X1
xU6140 n3611 n3703 n3702 VDD GND XOR2_X1
xU6141 n3704 n3705 n3611 VDD GND XOR2_X1
xU6142 n453 n3706 n3699 VDD GND XOR2_X1
xU6143 n3678 n3511 n3706 VDD GND XOR2_X1
xU6144 n3707 n3481 n3501 VDD GND XOR2_X1
xU6145 n735 Din_54 n3710 VDD GND XOR2_X1
xU6146 n3722 n3723 n3718 VDD GND XOR2_X1
xU6147 n471 n3724 n3723 VDD GND XOR2_X1
xU6148 n447 n3725 n3724 VDD GND XOR2_X1
xU6149 n290 n3726 n3722 VDD GND XOR2_X1
xU6150 n3727 n3728 n3726 VDD GND XOR2_X1
xU6151 n734 Din_53 n3731 VDD GND XOR2_X1
xU6152 n3744 n3745 n3740 VDD GND XOR2_X1
xU6153 n3746 n3747 n3745 VDD GND XOR2_X1
xU6154 n3748 n3749 n3747 VDD GND XOR2_X1
xU6155 n3583 n472 n3746 VDD GND XOR2_X1
xU6156 n3750 n3751 n3744 VDD GND XOR2_X1
xU6157 n3530 n3752 n3751 VDD GND XOR2_X1
xU6158 n3725 n3610 n3750 VDD GND XOR2_X1
xU6159 n733 Din_52 n3755 VDD GND XOR2_X1
xU6160 n3768 n3769 n3764 VDD GND XOR2_X1
xU6161 n3770 n3771 n3769 VDD GND XOR2_X1
xU6162 n3772 n3773 n3771 VDD GND XOR2_X1
xU6163 n3774 n3775 n3768 VDD GND XOR2_X1
xU6164 n3776 n3613 n3775 VDD GND XOR2_X1
xU6165 n3582 n297 n3613 VDD GND XOR2_X1
xU6166 n3777 n609 n3774 VDD GND XOR2_X1
xU6167 n732 Din_51 n3780 VDD GND XOR2_X1
xU6168 n3793 n3794 n3788 VDD GND XOR2_X1
xU6169 n3795 n298 n3793 VDD GND XOR2_X1
xU6170 n3796 n3797 n3789 VDD GND XOR2_X1
xU6171 n277 n3798 n3797 VDD GND XOR2_X1
xU6172 n3603 n3680 n3798 VDD GND XOR2_X1
xU6173 n3799 n3800 n3680 VDD GND XOR2_X1
xU6174 n3801 n3777 n3800 VDD GND XOR2_X1
xU6175 n3802 n3803 n3603 VDD GND XOR2_X1
xU6176 n3804 n3805 n3796 VDD GND XOR2_X1
xU6177 n3806 n3807 n3805 VDD GND XOR2_X1
xU6178 n3704 n3808 n3804 VDD GND XOR2_X1
xU6179 n731 Din_50 n3811 VDD GND XOR2_X1
xU6180 n3824 n3825 n3820 VDD GND XOR2_X1
xU6181 n3826 n3827 n3825 VDD GND XOR2_X1
xU6182 n3610 n3607 n3827 VDD GND XOR2_X1
xU6183 n612 n3828 n3607 VDD GND XOR2_X1
xU6184 n3772 n3829 n3824 VDD GND XOR2_X1
xU6185 n3656 n3830 n3829 VDD GND XOR2_X1
xU6186 n3831 n3832 n3656 VDD GND XOR2_X1
xU6187 n3583 n3833 n3832 VDD GND XOR2_X1
xU6188 n3834 n3835 n3831 VDD GND XOR2_X1
xU6189 n3509 n3531 n3835 VDD GND XOR2_X1
xU6190 n3836 n3658 n3772 VDD GND XOR2_X1
xU6191 n730 Din_49 n3839 VDD GND XOR2_X1
xU6192 n3852 n3853 n3848 VDD GND XOR2_X1
xU6193 n3854 n3855 n3853 VDD GND XOR2_X1
xU6194 n3856 n451 n3852 VDD GND XOR2_X1
xU6195 n729 Din_48 n3859 VDD GND XOR2_X1
xU6196 n3482 n3801 n3867 VDD GND XOR2_X1
xU6197 n3872 n3873 n3868 VDD GND XOR2_X1
xU6198 n3670 n3874 n3873 VDD GND XOR2_X1
xU6199 n3476 n3507 n3874 VDD GND XOR2_X1
xU6200 n3704 n3875 n3507 VDD GND XOR2_X1
xU6201 n3876 n3877 n3476 VDD GND XOR2_X1
xU6202 n3659 n3878 n3670 VDD GND XOR2_X1
xU6203 n3879 n3880 n3872 VDD GND XOR2_X1
xU6204 n728 Din_47 n3883 VDD GND XOR2_X1
xU6205 n3896 n3897 n3891 VDD GND XOR2_X1
xU6206 n603 n3898 n3897 VDD GND XOR2_X1
xU6207 n3481 n3698 n3898 VDD GND XOR2_X1
xU6208 n3899 n3900 n3896 VDD GND XOR2_X1
xU6209 n3901 n3880 n3900 VDD GND XOR2_X1
xU6210 n3902 n3903 n3880 VDD GND XOR2_X1
xU6211 n727 Din_46 n3906 VDD GND XOR2_X1
xU6212 n3918 n3919 n3914 VDD GND XOR2_X1
xU6213 n3920 n3921 n3919 VDD GND XOR2_X1
xU6214 n3504 n481 n3921 VDD GND XOR2_X1
xU6215 n3922 n3877 n3504 VDD GND XOR2_X1
xU6216 n3923 n3701 n3918 VDD GND XOR2_X1
xU6217 n478 n3557 n3923 VDD GND XOR2_X1
xU6218 n726 Din_45 n3926 VDD GND XOR2_X1
xU6219 n3938 n3939 n3934 VDD GND XOR2_X1
xU6220 n3940 n3941 n3939 VDD GND XOR2_X1
xU6221 n290 n3942 n3941 VDD GND XOR2_X1
xU6222 n3943 n3944 n3938 VDD GND XOR2_X1
xU6223 n3530 n3945 n3944 VDD GND XOR2_X1
xU6224 n3946 n3947 n3530 VDD GND XOR2_X1
xU6225 n454 n3948 n3947 VDD GND XOR2_X1
xU6226 n3949 n3950 n3946 VDD GND XOR2_X1
xU6227 n3951 n3952 n3949 VDD GND XOR2_X1
xU6228 n3836 n3953 n3943 VDD GND XOR2_X1
xU6229 n725 Din_44 n3956 VDD GND XOR2_X1
xU6230 n3968 n3969 n3964 VDD GND XOR2_X1
xU6231 n3970 n3971 n3969 VDD GND XOR2_X1
xU6232 n3770 n3972 n3971 VDD GND XOR2_X1
xU6233 n450 n3808 n3770 VDD GND XOR2_X1
xU6234 n3973 n608 n3970 VDD GND XOR2_X1
xU6235 n3974 n3975 n3968 VDD GND XOR2_X1
xU6236 n3976 n3704 n3975 VDD GND XOR2_X1
xU6237 n609 n3977 n3704 VDD GND XOR2_X1
xU6238 n3978 n612 n3974 VDD GND XOR2_X1
xU6239 n724 Din_43 n3981 VDD GND XOR2_X1
xU6240 n3994 n3995 n3989 VDD GND XOR2_X1
xU6241 n3801 n612 n3994 VDD GND XOR2_X1
xU6242 n3996 n3997 n3990 VDD GND XOR2_X1
xU6243 n3998 n3999 n3997 VDD GND XOR2_X1
xU6244 n3879 n3899 n3999 VDD GND XOR2_X1
xU6245 n3485 n3977 n3899 VDD GND XOR2_X1
xU6246 n3976 n3799 n3879 VDD GND XOR2_X1
xU6247 n3794 n4000 n3998 VDD GND XOR2_X1
xU6248 n3659 n4001 n3794 VDD GND XOR2_X1
xU6249 n4002 n4003 n3996 VDD GND XOR2_X1
xU6250 n4004 n3803 n4003 VDD GND XOR2_X1
xU6251 n473 n456 n4002 VDD GND XOR2_X1
xU6252 n723 Din_42 n4007 VDD GND XOR2_X1
xU6253 n4020 n3942 n4015 VDD GND XOR2_X1
xU6254 n4021 n4022 n4016 VDD GND XOR2_X1
xU6255 n4023 n4024 n4022 VDD GND XOR2_X1
xU6256 n3973 n3828 n4024 VDD GND XOR2_X1
xU6257 n3806 n3553 n3828 VDD GND XOR2_X1
xU6258 n452 n3877 n3553 VDD GND XOR2_X1
xU6259 n4004 n4025 n3877 VDD GND XOR2_X1
xU6260 n4026 n4027 n4021 VDD GND XOR2_X1
xU6261 n3819 n3854 n4027 VDD GND XOR2_X1
xU6262 n4028 n4029 n3854 VDD GND XOR2_X1
xU6263 n4030 n4031 n4029 VDD GND XOR2_X1
xU6264 n3836 n4032 n4031 VDD GND XOR2_X1
xU6265 n4033 n4034 n4028 VDD GND XOR2_X1
xU6266 n3678 n3725 n4034 VDD GND XOR2_X1
xU6267 n4035 n3749 n3819 VDD GND XOR2_X1
xU6268 n722 Din_41 n4038 VDD GND XOR2_X1
xU6269 n4051 n4052 n4047 VDD GND XOR2_X1
xU6270 n3847 n4053 n4052 VDD GND XOR2_X1
xU6271 n451 n3482 n4053 VDD GND XOR2_X1
xU6272 n3570 n4054 n3648 VDD GND XOR2_X1
xU6273 n3940 n4055 n4051 VDD GND XOR2_X1
xU6274 n481 n4026 n3940 VDD GND XOR2_X1
xU6275 n4056 n3801 n4026 VDD GND XOR2_X1
xU6276 n721 Din_40 n4059 VDD GND XOR2_X1
xU6277 n4056 n3679 n3479 VDD GND XOR2_X1
xU6278 n4071 n4072 n4067 VDD GND XOR2_X1
xU6279 n4073 n4074 n4072 VDD GND XOR2_X1
xU6280 n3802 n3855 n4074 VDD GND XOR2_X1
xU6281 n3610 n3878 n3855 VDD GND XOR2_X1
xU6282 n4075 n3585 n3878 VDD GND XOR2_X1
xU6283 n445 n3707 n3802 VDD GND XOR2_X1
xU6284 n4076 n4077 n4071 VDD GND XOR2_X1
xU6285 n3511 n3482 n4077 VDD GND XOR2_X1
xU6286 n4078 n3777 n3482 VDD GND XOR2_X1
xU6287 n455 n4079 n4076 VDD GND XOR2_X1
xU6288 n720 Din_39 n4082 VDD GND XOR2_X1
xU6289 n3977 n3511 n4090 VDD GND XOR2_X1
xU6290 n4095 n4096 n4091 VDD GND XOR2_X1
xU6291 n610 n4097 n4096 VDD GND XOR2_X1
xU6292 n4098 n3922 n4097 VDD GND XOR2_X1
xU6293 n4099 n4100 n3922 VDD GND XOR2_X1
xU6294 n4101 n3875 n3895 VDD GND XOR2_X1
xU6295 n4102 n4103 n4095 VDD GND XOR2_X1
xU6296 n3485 n445 n4103 VDD GND XOR2_X1
xU6297 n4104 n3950 n4004 VDD GND XOR2_X1
xU6298 n4105 n4106 n3950 VDD GND XOR2_X1
xU6299 n3698 n4079 n4102 VDD GND XOR2_X1
xU6300 n719 Din_38 n4109 VDD GND XOR2_X1
xU6301 n4121 n3901 n4098 VDD GND XOR2_X1
xU6302 n4122 n3945 n3901 VDD GND XOR2_X1
xU6303 n4123 n4124 n3945 VDD GND XOR2_X1
xU6304 n4125 n4126 n4117 VDD GND XOR2_X1
xU6305 n269 n4127 n4126 VDD GND XOR2_X1
xU6306 n450 n472 n4127 VDD GND XOR2_X1
xU6307 n3558 n3803 n3570 VDD GND XOR2_X1
xU6308 n3876 n4128 n3803 VDD GND XOR2_X1
xU6309 n4075 n3506 n3701 VDD GND XOR2_X1
xU6310 n4129 n3554 n3506 VDD GND XOR2_X1
xU6311 n4130 n4131 n3554 VDD GND XOR2_X1
xU6312 n3528 n4132 n4125 VDD GND XOR2_X1
xU6313 n4104 n4133 n4132 VDD GND XOR2_X1
xU6314 n4078 n3703 n3528 VDD GND XOR2_X1
xU6315 n4134 n3752 n3703 VDD GND XOR2_X1
xU6316 n4135 n4136 n3752 VDD GND XOR2_X1
xU6317 n718 Din_37 n4139 VDD GND XOR2_X1
xU6318 n4152 n4153 n4147 VDD GND XOR2_X1
xU6319 n473 n3953 n4153 VDD GND XOR2_X1
xU6320 n3920 n4154 n3953 VDD GND XOR2_X1
xU6321 n4155 n4156 n3920 VDD GND XOR2_X1
xU6322 n4157 n4158 n4156 VDD GND XOR2_X1
xU6323 n485 n4161 n4159 VDD GND XOR2_X1
xU6324 n4162 n4163 n4152 VDD GND XOR2_X1
xU6325 n4164 n4165 n4162 VDD GND XOR2_X1
xU6326 n4166 n4167 n4148 VDD GND XOR2_X1
xU6327 n4168 n4169 n4167 VDD GND XOR2_X1
xU6328 n3557 n3948 n4169 VDD GND XOR2_X1
xU6329 n4133 n4170 n3948 VDD GND XOR2_X1
xU6330 n4171 n4172 n4133 VDD GND XOR2_X1
xU6331 n4173 n4174 n4172 VDD GND XOR2_X1
xU6332 Dout_E_57 n4177 n4175 VDD GND XOR2_X1
xU6333 n4178 n4179 n3557 VDD GND XOR2_X1
xU6334 n3808 n3748 n4179 VDD GND XOR2_X1
xU6335 n3727 n4180 n3748 VDD GND XOR2_X1
xU6336 n4181 n4182 n3727 VDD GND XOR2_X1
xU6337 n4183 n4184 n4182 VDD GND XOR2_X1
xU6338 n618 n4187 n4185 VDD GND XOR2_X1
xU6339 n4188 n4189 n4178 VDD GND XOR2_X1
xU6340 n4190 n4191 n4188 VDD GND XOR2_X1
xU6341 n4104 n4100 n4168 VDD GND XOR2_X1
xU6342 n4192 n4193 n4100 VDD GND XOR2_X1
xU6343 n4194 n4195 n4166 VDD GND XOR2_X1
xU6344 n3973 n3826 n4195 VDD GND XOR2_X1
xU6345 n290 n3799 n4194 VDD GND XOR2_X1
xU6346 n4196 n4197 n3739 VDD GND XOR2_X1
xU6347 n3552 n3582 n4197 VDD GND XOR2_X1
xU6348 n3533 n4198 n3552 VDD GND XOR2_X1
xU6349 n4199 n4200 n3533 VDD GND XOR2_X1
xU6350 n4201 n4202 n4200 VDD GND XOR2_X1
xU6351 Dout_E_17 n4205 n4203 VDD GND XOR2_X1
xU6352 n4206 n4207 n4196 VDD GND XOR2_X1
xU6353 n4208 n4209 n4206 VDD GND XOR2_X1
xU6354 n717 Din_36 n4212 VDD GND XOR2_X1
xU6355 n4224 n4225 n4220 VDD GND XOR2_X1
xU6356 n4073 n4226 n4225 VDD GND XOR2_X1
xU6357 n3806 n3972 n4226 VDD GND XOR2_X1
xU6358 n262 n4227 n3972 VDD GND XOR2_X1
xU6359 n456 n477 n3806 VDD GND XOR2_X1
xU6360 n3876 n3977 n4073 VDD GND XOR2_X1
xU6361 n4228 n4229 n4224 VDD GND XOR2_X1
xU6362 n4230 n3580 n4229 VDD GND XOR2_X1
xU6363 n602 n4025 n3580 VDD GND XOR2_X1
xU6364 n3558 n3707 n4228 VDD GND XOR2_X1
xU6365 n716 Din_35 n4233 VDD GND XOR2_X1
xU6366 n4246 n3614 n4241 VDD GND XOR2_X1
xU6367 n4056 n3807 n3614 VDD GND XOR2_X1
xU6368 n480 n4247 n3807 VDD GND XOR2_X1
xU6369 n3977 n477 n4246 VDD GND XOR2_X1
xU6370 n4248 n4249 n3977 VDD GND XOR2_X1
xU6371 n4250 n4157 n4249 VDD GND XOR2_X1
xU6372 n485 n4253 n4251 VDD GND XOR2_X1
xU6373 n470 n4256 n4242 VDD GND XOR2_X1
xU6374 n4257 n4258 n4256 VDD GND XOR2_X1
xU6375 n4259 n4260 n4258 VDD GND XOR2_X1
xU6376 n4001 n3995 n4260 VDD GND XOR2_X1
xU6377 n3682 n3609 n3995 VDD GND XOR2_X1
xU6378 n609 n3705 n3682 VDD GND XOR2_X1
xU6379 n4261 n4262 n4101 VDD GND XOR2_X1
xU6380 n4263 n4183 n4262 VDD GND XOR2_X1
xU6381 n618 n4266 n4264 VDD GND XOR2_X1
xU6382 n285 n4269 n4001 VDD GND XOR2_X1
xU6383 n3876 n3773 n4259 VDD GND XOR2_X1
xU6384 n4099 n4170 n3876 VDD GND XOR2_X1
xU6385 n4274 n4275 n4257 VDD GND XOR2_X1
xU6386 n454 n3610 n4275 VDD GND XOR2_X1
xU6387 n3659 n3801 n3610 VDD GND XOR2_X1
xU6388 n3481 n4079 n4025 VDD GND XOR2_X1
xU6389 n3485 n455 n4274 VDD GND XOR2_X1
xU6390 n297 n3707 n3485 VDD GND XOR2_X1
xU6391 n4280 n4281 n3707 VDD GND XOR2_X1
xU6392 n4282 n4173 n4281 VDD GND XOR2_X1
xU6393 n460 n4285 n4283 VDD GND XOR2_X1
xU6394 n4288 n4289 n3795 VDD GND XOR2_X1
xU6395 n4290 n4201 n4289 VDD GND XOR2_X1
xU6396 n303 n304 n4291 VDD GND XOR2_X1
xU6397 n715 Din_34 n4297 VDD GND XOR2_X1
xU6398 n3978 n3826 n3637 VDD GND XOR2_X1
xU6399 n4121 n4230 n3826 VDD GND XOR2_X1
xU6400 n4310 n4311 n4305 VDD GND XOR2_X1
xU6401 n4312 n4313 n4311 VDD GND XOR2_X1
xU6402 n4054 n3632 n4313 VDD GND XOR2_X1
xU6403 n3558 n4000 n3632 VDD GND XOR2_X1
xU6404 n3773 n3942 n4000 VDD GND XOR2_X1
xU6405 n4078 n608 n3942 VDD GND XOR2_X1
xU6406 n3808 n3705 n4078 VDD GND XOR2_X1
xU6407 n3725 n4189 n3705 VDD GND XOR2_X1
xU6408 n4033 n4314 n4189 VDD GND XOR2_X1
xU6409 Dout_E_105 n4317 n4316 VDD GND XOR2_X1
xU6410 n3875 n3678 n3808 VDD GND XOR2_X1
xU6411 n298 n612 n3773 VDD GND XOR2_X1
xU6412 n4322 n4323 n4054 VDD GND XOR2_X1
xU6413 n3481 n4106 n4322 VDD GND XOR2_X1
xU6414 n3586 n481 n4312 VDD GND XOR2_X1
xU6415 n4055 n4327 n4310 VDD GND XOR2_X1
xU6416 n3799 n3749 n4327 VDD GND XOR2_X1
xU6417 n4075 n3658 n3749 VDD GND XOR2_X1
xU6418 n3582 n3510 n4075 VDD GND XOR2_X1
xU6419 n3531 n4207 n3510 VDD GND XOR2_X1
xU6420 n3834 n4328 n4207 VDD GND XOR2_X1
xU6421 Dout_E_17 n4332 n4330 VDD GND XOR2_X1
xU6422 n3698 n3509 n3582 VDD GND XOR2_X1
xU6423 n4335 n4336 n4055 VDD GND XOR2_X1
xU6424 n3973 n4337 n4336 VDD GND XOR2_X1
xU6425 n4338 n4230 n4335 VDD GND XOR2_X1
xU6426 n4339 n3902 n4338 VDD GND XOR2_X1
xU6427 n714 Din_33 n4342 VDD GND XOR2_X1
xU6428 n3776 n4023 n3856 VDD GND XOR2_X1
xU6429 n4354 n4337 n4023 VDD GND XOR2_X1
xU6430 n4248 n4155 n4337 VDD GND XOR2_X1
xU6431 n3511 n4358 n4354 VDD GND XOR2_X1
xU6432 n4247 n3973 n3776 VDD GND XOR2_X1
xU6433 n4123 n4164 n3973 VDD GND XOR2_X1
xU6434 n3976 n4230 n4247 VDD GND XOR2_X1
xU6435 n4124 n4165 n4230 VDD GND XOR2_X1
xU6436 n4363 n4364 n4350 VDD GND XOR2_X1
xU6437 n257 n4365 n4364 VDD GND XOR2_X1
xU6438 n601 n3799 n4365 VDD GND XOR2_X1
xU6439 n455 n4056 n3799 VDD GND XOR2_X1
xU6440 n4176 n4270 n4324 VDD GND XOR2_X1
xU6441 n4369 n4370 n4270 VDD GND XOR2_X1
xU6442 n602 n3830 n4046 VDD GND XOR2_X1
xU6443 n4373 n4030 n3830 VDD GND XOR2_X1
xU6444 n4261 n4181 n4030 VDD GND XOR2_X1
xU6445 n3875 n4314 n4373 VDD GND XOR2_X1
xU6446 n4186 n613 n4276 VDD GND XOR2_X1
xU6447 n3836 n3609 n3728 VDD GND XOR2_X1
xU6448 n3777 n4032 n3609 VDD GND XOR2_X1
xU6449 n4136 n4191 n4032 VDD GND XOR2_X1
xU6450 n4134 n4180 n3777 VDD GND XOR2_X1
xU6451 n4380 n4381 n4375 VDD GND XOR2_X1
xU6452 n4267 n4318 n4374 VDD GND XOR2_X1
xU6453 n4383 n4380 n4318 VDD GND XOR2_X1
xU6454 n4135 n4190 n3836 VDD GND XOR2_X1
xU6455 n4389 n4390 n4384 VDD GND XOR2_X1
xU6456 n4391 n4392 n4390 VDD GND XOR2_X1
xU6457 n4265 n611 n4315 VDD GND XOR2_X1
xU6458 n4383 n4381 n4394 VDD GND XOR2_X1
xU6459 n4398 n4399 n4389 VDD GND XOR2_X1
xU6460 n4400 n4266 n4399 VDD GND XOR2_X1
xU6461 n4401 n4402 n4395 VDD GND XOR2_X1
xU6462 n4391 n4403 n4402 VDD GND XOR2_X1
xU6463 n4406 n4407 n4405 VDD GND XOR2_X1
xU6464 n4408 n4409 n4407 VDD GND XOR2_X1
xU6465 n4410 n4411 n4404 VDD GND XOR2_X1
xU6466 n4187 n4409 n4411 VDD GND XOR2_X1
xU6467 n4412 n4413 n4409 VDD GND XOR2_X1
xU6468 n4406 n4414 n4401 VDD GND XOR2_X1
xU6469 n4415 n4410 n4414 VDD GND XOR2_X1
xU6470 n4416 n4417 n4410 VDD GND XOR2_X1
xU6471 n4418 n4419 n4406 VDD GND XOR2_X1
xU6472 n4388 n4420 n4397 VDD GND XOR2_X1
xU6473 n4403 n4392 n4420 VDD GND XOR2_X1
xU6474 n619 n4421 n4396 VDD GND XOR2_X1
xU6475 n4398 n4422 n4421 VDD GND XOR2_X1
xU6476 n4418 n4423 n4398 VDD GND XOR2_X1
xU6477 n617 n4266 n4424 VDD GND XOR2_X1
xU6478 n4317 Dout_E_104 n4393 VDD GND XOR2_X1
xU6479 n4408 n620 n4187 VDD GND XOR2_X1
xU6480 n4268 n4426 n4425 VDD GND XOR2_X1
xU6481 n4422 n4400 n4426 VDD GND XOR2_X1
xU6482 n4417 n4427 n4400 VDD GND XOR2_X1
xU6483 Dout_E_105 n4429 n4428 VDD GND XOR2_X1
xU6484 n4317 n4429 n4378 VDD GND XOR2_X1
xU6485 Dout_E_109 n4430 n4317 VDD GND XOR2_X1
xU6486 n4431 n4413 n4422 VDD GND XOR2_X1
xU6487 Dout_E_107 n624 n4432 VDD GND XOR2_X1
xU6488 Dout_E_109 Dout_E_111 n4268 VDD GND XOR2_X1
xU6489 n4434 n4435 n4385 VDD GND XOR2_X1
xU6490 n620 n4436 n4434 VDD GND XOR2_X1
xU6491 n616 n4437 n4433 VDD GND XOR2_X1
xU6492 n4435 n4266 n4437 VDD GND XOR2_X1
xU6493 n4438 n4430 n4266 VDD GND XOR2_X1
xU6494 n4412 n4431 n4435 VDD GND XOR2_X1
xU6495 n4440 n4441 n4439 VDD GND XOR2_X1
xU6496 Dout_E_111 Dout_E_110 n4441 VDD GND XOR2_X1
xU6497 Dout_E_110 n4320 n4386 VDD GND XOR2_X1
xU6498 Dout_E_109 n4440 n4320 VDD GND XOR2_X1
xU6499 n621 n618 n4440 VDD GND XOR2_X1
xU6500 Dout_E_108 n4443 n4442 VDD GND XOR2_X1
xU6501 n4445 n4446 n4388 VDD GND XOR2_X1
xU6502 n4438 n4444 n4446 VDD GND XOR2_X1
xU6503 n4416 n4427 n4444 VDD GND XOR2_X1
xU6504 Dout_E_105 n4447 n4379 VDD GND XOR2_X1
xU6505 n623 n4443 n4319 VDD GND XOR2_X1
xU6506 Dout_E_105 n4430 n4443 VDD GND XOR2_X1
xU6507 n628 n4415 n4430 VDD GND XOR2_X1
xU6508 n621 Dout_E_107 n4415 VDD GND XOR2_X1
xU6509 n626 n624 n4408 VDD GND XOR2_X1
xU6510 n625 Dout_E_110 n4438 VDD GND XOR2_X1
xU6511 n628 n4436 n4445 VDD GND XOR2_X1
xU6512 n4423 n4419 n4436 VDD GND XOR2_X1
xU6513 Dout_E_106 n4451 n4450 VDD GND XOR2_X1
xU6514 Dout_E_107 n4451 n4382 VDD GND XOR2_X1
xU6515 n625 n628 n4451 VDD GND XOR2_X1
xU6516 n4453 n4447 n4277 VDD GND XOR2_X1
xU6517 n617 n625 n4447 VDD GND XOR2_X1
xU6518 n621 n626 n4453 VDD GND XOR2_X1
xU6519 Dout_E_107 n4429 n4452 VDD GND XOR2_X1
xU6520 n617 n627 n4429 VDD GND XOR2_X1
xU6521 n3763 n3634 n3847 VDD GND XOR2_X1
xU6522 n4454 n3833 n3634 VDD GND XOR2_X1
xU6523 n4288 n4199 n3833 VDD GND XOR2_X1
xU6524 n3698 n4328 n4454 VDD GND XOR2_X1
xU6525 n4204 n4456 n4278 VDD GND XOR2_X1
xU6526 n3583 n4269 n3763 VDD GND XOR2_X1
xU6527 n3585 n3658 n4269 VDD GND XOR2_X1
xU6528 n4131 n4209 n3658 VDD GND XOR2_X1
xU6529 n4129 n4198 n3585 VDD GND XOR2_X1
xU6530 n4461 n4462 n4456 VDD GND XOR2_X1
xU6531 n4293 n4333 n4455 VDD GND XOR2_X1
xU6532 n4462 n4464 n4333 VDD GND XOR2_X1
xU6533 n4130 n4208 n3583 VDD GND XOR2_X1
xU6534 n4470 n4471 n4466 VDD GND XOR2_X1
xU6535 n4472 n4473 n4471 VDD GND XOR2_X1
xU6536 n4292 n4331 n4329 VDD GND XOR2_X1
xU6537 n4461 n4464 n4331 VDD GND XOR2_X1
xU6538 n299 n4479 n4470 VDD GND XOR2_X1
xU6539 n4480 n304 n4479 VDD GND XOR2_X1
xU6540 n4482 n4483 n4478 VDD GND XOR2_X1
xU6541 n4472 n4484 n4483 VDD GND XOR2_X1
xU6542 n4486 n4487 n4476 VDD GND XOR2_X1
xU6543 n4488 n4489 n4487 VDD GND XOR2_X1
xU6544 n4490 n4491 n4486 VDD GND XOR2_X1
xU6545 n4492 n4493 n4485 VDD GND XOR2_X1
xU6546 n4491 n4494 n4493 VDD GND XOR2_X1
xU6547 n4494 n4495 n4482 VDD GND XOR2_X1
xU6548 n4496 n4488 n4495 VDD GND XOR2_X1
xU6549 n4497 n4498 n4488 VDD GND XOR2_X1
xU6550 n302 n4499 n4494 VDD GND XOR2_X1
xU6551 n4469 n4501 n4475 VDD GND XOR2_X1
xU6552 n4484 n4473 n4501 VDD GND XOR2_X1
xU6553 n4492 n4503 n4477 VDD GND XOR2_X1
xU6554 n4504 n4481 n4503 VDD GND XOR2_X1
xU6555 n4497 n4505 n4481 VDD GND XOR2_X1
xU6556 n301 n304 n4506 VDD GND XOR2_X1
xU6557 n4332 Dout_E_16 n4474 VDD GND XOR2_X1
xU6558 n4205 n4490 n4492 VDD GND XOR2_X1
xU6559 n308 n305 n4205 VDD GND XOR2_X1
xU6560 n4508 n4509 n4502 VDD GND XOR2_X1
xU6561 n4294 n4480 n4509 VDD GND XOR2_X1
xU6562 n4499 n4510 n4480 VDD GND XOR2_X1
xU6563 Dout_E_17 n4512 n4511 VDD GND XOR2_X1
xU6564 n4332 n4512 n4459 VDD GND XOR2_X1
xU6565 Dout_E_21 n4513 n4332 VDD GND XOR2_X1
xU6566 Dout_E_21 Dout_E_23 n4294 VDD GND XOR2_X1
xU6567 n4504 n4490 n4508 VDD GND XOR2_X1
xU6568 Dout_E_19 n4515 n4514 VDD GND XOR2_X1
xU6569 Dout_E_17 n4516 n4321 VDD GND XOR2_X1
xU6570 n4518 n4519 n4465 VDD GND XOR2_X1
xU6571 n305 n4520 n4519 VDD GND XOR2_X1
xU6572 n4521 n4522 n4517 VDD GND XOR2_X1
xU6573 n4507 n4520 n4522 VDD GND XOR2_X1
xU6574 n4491 n4504 n4520 VDD GND XOR2_X1
xU6575 n4524 n4525 n4523 VDD GND XOR2_X1
xU6576 n4516 n4525 n4467 VDD GND XOR2_X1
xU6577 n311 n303 n4525 VDD GND XOR2_X1
xU6578 Dout_E_20 n4527 n4526 VDD GND XOR2_X1
xU6579 n4515 n4513 n4507 VDD GND XOR2_X1
xU6580 n4528 n4529 n4469 VDD GND XOR2_X1
xU6581 n4518 n4521 n4529 VDD GND XOR2_X1
xU6582 n4500 n4510 n4521 VDD GND XOR2_X1
xU6583 Dout_E_17 n4530 n4460 VDD GND XOR2_X1
xU6584 n308 n4527 n4334 VDD GND XOR2_X1
xU6585 Dout_E_17 n4513 n4527 VDD GND XOR2_X1
xU6586 n312 n4496 n4513 VDD GND XOR2_X1
xU6587 n306 Dout_E_19 n4496 VDD GND XOR2_X1
xU6588 n310 n4515 n4489 VDD GND XOR2_X1
xU6589 n4505 n4498 n4518 VDD GND XOR2_X1
xU6590 Dout_E_19 n4534 n4463 VDD GND XOR2_X1
xU6591 Dout_E_23 Dout_E_20 n4534 VDD GND XOR2_X1
xU6592 Dout_E_20 n4524 n4533 VDD GND XOR2_X1
xU6593 n306 n312 n4524 VDD GND XOR2_X1
xU6594 n4516 n4530 n4279 VDD GND XOR2_X1
xU6595 n301 n309 n4530 VDD GND XOR2_X1
xU6596 Dout_E_18 Dout_E_21 n4516 VDD GND XOR2_X1
xU6597 Dout_E_19 n4512 n4535 VDD GND XOR2_X1
xU6598 n301 n311 n4512 VDD GND XOR2_X1
xU6599 Dout_E_23 n4515 n4528 VDD GND XOR2_X1
xU6600 Dout_E_20 Dout_E_22 n4515 VDD GND XOR2_X1
xU6601 n3636 n4536 n4363 VDD GND XOR2_X1
xU6602 n3679 n3558 n4536 VDD GND XOR2_X1
xU6603 n4192 n3951 n3558 VDD GND XOR2_X1
xU6604 n4121 n3976 n3679 VDD GND XOR2_X1
xU6605 n4122 n4154 n3976 VDD GND XOR2_X1
xU6606 n4254 n4355 n4357 VDD GND XOR2_X1
xU6607 n473 n480 n4121 VDD GND XOR2_X1
xU6608 n4325 n4163 n3903 VDD GND XOR2_X1
xU6609 n4339 n4358 n4163 VDD GND XOR2_X1
xU6610 n4252 n482 n4360 VDD GND XOR2_X1
xU6611 n4551 n4552 n4550 VDD GND XOR2_X1
xU6612 Dout_E_65 n4356 n4549 VDD GND XOR2_X1
xU6613 n3511 n3902 n4227 VDD GND XOR2_X1
xU6614 n4551 n4554 n4355 VDD GND XOR2_X1
xU6615 n4556 n4557 n4547 VDD GND XOR2_X1
xU6616 n4558 n4559 n4557 VDD GND XOR2_X1
xU6617 n4160 n479 n4366 VDD GND XOR2_X1
xU6618 n4554 n4552 n4544 VDD GND XOR2_X1
xU6619 n4565 n4548 n4560 VDD GND XOR2_X1
xU6620 n4566 n4567 n4548 VDD GND XOR2_X1
xU6621 n488 n4568 n4567 VDD GND XOR2_X1
xU6622 n4572 n4573 n4563 VDD GND XOR2_X1
xU6623 n4569 n4574 n4572 VDD GND XOR2_X1
xU6624 n4575 n4576 n4571 VDD GND XOR2_X1
xU6625 n486 n4577 n4575 VDD GND XOR2_X1
xU6626 n4564 n4578 n4562 VDD GND XOR2_X1
xU6627 n4570 n4559 n4578 VDD GND XOR2_X1
xU6628 n4161 n4580 n4561 VDD GND XOR2_X1
xU6629 n4574 n4581 n4580 VDD GND XOR2_X1
xU6630 n4582 n4583 n4574 VDD GND XOR2_X1
xU6631 n4577 n4584 n4579 VDD GND XOR2_X1
xU6632 n4255 n4585 n4584 VDD GND XOR2_X1
xU6633 Dout_E_69 Dout_E_71 n4255 VDD GND XOR2_X1
xU6634 n4582 n4586 n4577 VDD GND XOR2_X1
xU6635 n4588 n4589 n4587 VDD GND XOR2_X1
xU6636 Dout_E_71 Dout_E_66 n4589 VDD GND XOR2_X1
xU6637 n4588 n4590 n4359 VDD GND XOR2_X1
xU6638 Dout_E_70 Dout_E_65 n4588 VDD GND XOR2_X1
xU6639 n4545 n4592 n4555 VDD GND XOR2_X1
xU6640 n4573 n4581 n4592 VDD GND XOR2_X1
xU6641 n4593 n4594 n4581 VDD GND XOR2_X1
xU6642 n4595 n4596 n4573 VDD GND XOR2_X1
xU6643 n484 n4597 n4591 VDD GND XOR2_X1
xU6644 n4161 n4585 n4597 VDD GND XOR2_X1
xU6645 n4598 n4594 n4585 VDD GND XOR2_X1
xU6646 Dout_E_67 n491 n4599 VDD GND XOR2_X1
xU6647 Dout_E_65 n4590 n4309 VDD GND XOR2_X1
xU6648 n4545 n4569 n4161 VDD GND XOR2_X1
xU6649 n4600 n4595 n4576 VDD GND XOR2_X1
xU6650 Dout_E_68 n4602 n4601 VDD GND XOR2_X1
xU6651 n4568 n4603 n4564 VDD GND XOR2_X1
xU6652 n4604 n4253 n4603 VDD GND XOR2_X1
xU6653 n4593 n4598 n4568 VDD GND XOR2_X1
xU6654 Dout_E_65 n4606 n4605 VDD GND XOR2_X1
xU6655 n4356 n4606 n4362 VDD GND XOR2_X1
xU6656 n483 n4253 n4607 VDD GND XOR2_X1
xU6657 n4608 n4609 n4253 VDD GND XOR2_X1
xU6658 n4356 Dout_E_64 n4361 VDD GND XOR2_X1
xU6659 Dout_E_69 n4609 n4356 VDD GND XOR2_X1
xU6660 n4610 n4611 n4556 VDD GND XOR2_X1
xU6661 n4608 n4566 n4611 VDD GND XOR2_X1
xU6662 n4600 n4596 n4566 VDD GND XOR2_X1
xU6663 Dout_E_66 n4613 n4612 VDD GND XOR2_X1
xU6664 Dout_E_67 n4613 n4541 VDD GND XOR2_X1
xU6665 n492 n495 n4613 VDD GND XOR2_X1
xU6666 n4545 n4602 n4553 VDD GND XOR2_X1
xU6667 Dout_E_65 n4609 n4602 VDD GND XOR2_X1
xU6668 n495 n4569 n4609 VDD GND XOR2_X1
xU6669 n489 Dout_E_67 n4569 VDD GND XOR2_X1
xU6670 Dout_E_69 n491 n4545 VDD GND XOR2_X1
xU6671 n492 Dout_E_70 n4608 VDD GND XOR2_X1
xU6672 Dout_E_71 n4604 n4610 VDD GND XOR2_X1
xU6673 n4583 n4586 n4604 VDD GND XOR2_X1
xU6674 Dout_E_65 n4616 n4540 VDD GND XOR2_X1
xU6675 n4590 n4616 n4367 VDD GND XOR2_X1
xU6676 n483 n492 n4616 VDD GND XOR2_X1
xU6677 Dout_E_66 Dout_E_69 n4590 VDD GND XOR2_X1
xU6678 Dout_E_67 n4606 n4617 VDD GND XOR2_X1
xU6679 n483 n494 n4606 VDD GND XOR2_X1
xU6680 n4618 n4619 n3636 VDD GND XOR2_X1
xU6681 n452 n4323 n4619 VDD GND XOR2_X1
xU6682 n4280 n4171 n4323 VDD GND XOR2_X1
xU6683 n4286 n4620 n4272 VDD GND XOR2_X1
xU6684 n4193 n3952 n4128 VDD GND XOR2_X1
xU6685 n4105 n4626 n4618 VDD GND XOR2_X1
xU6686 n4079 n4104 n4626 VDD GND XOR2_X1
xU6687 Dout_E_57 n4621 n4627 VDD GND XOR2_X1
xU6688 n4370 n4629 n4620 VDD GND XOR2_X1
xU6689 n4632 n4633 n4631 VDD GND XOR2_X1
xU6690 n4634 n4635 n4633 VDD GND XOR2_X1
xU6691 n4284 n4624 n4538 VDD GND XOR2_X1
xU6692 n4369 n4629 n4624 VDD GND XOR2_X1
xU6693 n4641 n4642 n4632 VDD GND XOR2_X1
xU6694 n4643 n4285 n4642 VDD GND XOR2_X1
xU6695 n4644 n4645 n4639 VDD GND XOR2_X1
xU6696 n4634 n4646 n4645 VDD GND XOR2_X1
xU6697 n4648 n4649 n4638 VDD GND XOR2_X1
xU6698 n4636 n4650 n4649 VDD GND XOR2_X1
xU6699 n4651 n4652 n4648 VDD GND XOR2_X1
xU6700 n4653 n4654 n4647 VDD GND XOR2_X1
xU6701 n4652 n4655 n4654 VDD GND XOR2_X1
xU6702 n4655 n4656 n4644 VDD GND XOR2_X1
xU6703 n4657 n4650 n4656 VDD GND XOR2_X1
xU6704 n4658 n4659 n4650 VDD GND XOR2_X1
xU6705 n4660 n4661 n4655 VDD GND XOR2_X1
xU6706 n4623 n4662 n4637 VDD GND XOR2_X1
xU6707 n4646 n4635 n4662 VDD GND XOR2_X1
xU6708 n4653 n4664 n4640 VDD GND XOR2_X1
xU6709 n4665 n4641 n4664 VDD GND XOR2_X1
xU6710 n4658 n4666 n4641 VDD GND XOR2_X1
xU6711 n459 n4285 n4667 VDD GND XOR2_X1
xU6712 n4621 Dout_E_56 n4539 VDD GND XOR2_X1
xU6713 n4651 n4177 n4653 VDD GND XOR2_X1
xU6714 n4636 n461 n4177 VDD GND XOR2_X1
xU6715 n4668 n4669 n4663 VDD GND XOR2_X1
xU6716 n4287 n4643 n4669 VDD GND XOR2_X1
xU6717 n4661 n4670 n4643 VDD GND XOR2_X1
xU6718 Dout_E_57 n4672 n4671 VDD GND XOR2_X1
xU6719 n4621 n4672 n4625 VDD GND XOR2_X1
xU6720 Dout_E_61 n4673 n4621 VDD GND XOR2_X1
xU6721 Dout_E_61 Dout_E_63 n4287 VDD GND XOR2_X1
xU6722 n4651 n4665 n4668 VDD GND XOR2_X1
xU6723 Dout_E_59 n464 n4674 VDD GND XOR2_X1
xU6724 n4676 n4677 n4630 VDD GND XOR2_X1
xU6725 n4657 n4678 n4677 VDD GND XOR2_X1
xU6726 n4679 n4680 n4675 VDD GND XOR2_X1
xU6727 n4285 n4678 n4680 VDD GND XOR2_X1
xU6728 n4652 n4665 n4678 VDD GND XOR2_X1
xU6729 n4682 n4683 n4681 VDD GND XOR2_X1
xU6730 Dout_E_63 Dout_E_62 n4683 VDD GND XOR2_X1
xU6731 Dout_E_62 n4326 n4537 VDD GND XOR2_X1
xU6732 Dout_E_61 n4682 n4326 VDD GND XOR2_X1
xU6733 n462 n460 n4682 VDD GND XOR2_X1
xU6734 Dout_E_60 n4685 n4684 VDD GND XOR2_X1
xU6735 n4686 n4673 n4285 VDD GND XOR2_X1
xU6736 n4687 n4688 n4623 VDD GND XOR2_X1
xU6737 n4679 n4676 n4688 VDD GND XOR2_X1
xU6738 n4666 n4659 n4676 VDD GND XOR2_X1
xU6739 Dout_E_58 n4690 n4689 VDD GND XOR2_X1
xU6740 Dout_E_59 n4690 n4273 VDD GND XOR2_X1
xU6741 n465 n468 n4690 VDD GND XOR2_X1
xU6742 n4692 n4693 n4368 VDD GND XOR2_X1
xU6743 n462 n466 n4692 VDD GND XOR2_X1
xU6744 Dout_E_59 n4672 n4691 VDD GND XOR2_X1
xU6745 n459 n467 n4672 VDD GND XOR2_X1
xU6746 n4660 n4670 n4679 VDD GND XOR2_X1
xU6747 Dout_E_57 n4693 n4271 VDD GND XOR2_X1
xU6748 n459 n465 n4693 VDD GND XOR2_X1
xU6749 n4636 n4685 n4628 VDD GND XOR2_X1
xU6750 Dout_E_57 n4673 n4685 VDD GND XOR2_X1
xU6751 n468 n4657 n4673 VDD GND XOR2_X1
xU6752 n462 Dout_E_59 n4657 VDD GND XOR2_X1
xU6753 Dout_E_61 n464 n4636 VDD GND XOR2_X1
xU6754 n468 n4686 n4687 VDD GND XOR2_X1
xU6755 n465 Dout_E_62 n4686 VDD GND XOR2_X1
xU6756 n713 Din_32 n4698 VDD GND XOR2_X1
xU6757 n4711 n4712 n4706 VDD GND XOR2_X1
xU6758 n4713 n4714 n4707 VDD GND XOR2_X1
xU6759 n4715 n4716 n4714 VDD GND XOR2_X1
xU6760 n4717 n4718 n4716 VDD GND XOR2_X1
xU6761 n4719 n4720 n4715 VDD GND XOR2_X1
xU6762 n4721 n4722 n4713 VDD GND XOR2_X1
xU6763 n378 n4723 n4722 VDD GND XOR2_X1
xU6764 n4724 n4725 n4721 VDD GND XOR2_X1
xU6765 n712 Din_31 n4728 VDD GND XOR2_X1
xU6766 n352 n4719 n4736 VDD GND XOR2_X1
xU6767 n4741 n4742 n4737 VDD GND XOR2_X1
xU6768 n4743 n4744 n4742 VDD GND XOR2_X1
xU6769 n4745 n4746 n4744 VDD GND XOR2_X1
xU6770 n4747 n4748 n4741 VDD GND XOR2_X1
xU6771 n382 n4749 n4748 VDD GND XOR2_X1
xU6772 n4750 n4717 n4747 VDD GND XOR2_X1
xU6773 n711 Din_30 n4753 VDD GND XOR2_X1
xU6774 n4765 n4766 n4761 VDD GND XOR2_X1
xU6775 n374 n4767 n4766 VDD GND XOR2_X1
xU6776 n4768 n639 n4767 VDD GND XOR2_X1
xU6777 n499 n4769 n4765 VDD GND XOR2_X1
xU6778 n4770 n4771 n4769 VDD GND XOR2_X1
xU6779 n710 Din_29 n4774 VDD GND XOR2_X1
xU6780 n4786 n4787 n4782 VDD GND XOR2_X1
xU6781 n4788 n4789 n4787 VDD GND XOR2_X1
xU6782 n4790 n4791 n4789 VDD GND XOR2_X1
xU6783 n4792 n4770 n4788 VDD GND XOR2_X1
xU6784 n4793 n4794 n4786 VDD GND XOR2_X1
xU6785 n4795 n504 n4794 VDD GND XOR2_X1
xU6786 n4796 n356 n4793 VDD GND XOR2_X1
xU6787 n709 Din_28 n4799 VDD GND XOR2_X1
xU6788 n4812 n4813 n4807 VDD GND XOR2_X1
xU6789 n4814 n4815 n4813 VDD GND XOR2_X1
xU6790 n4816 n4817 n4815 VDD GND XOR2_X1
xU6791 n4818 n4819 n4812 VDD GND XOR2_X1
xU6792 n4724 n4820 n4818 VDD GND XOR2_X1
xU6793 n4821 n4822 n4724 VDD GND XOR2_X1
xU6794 n708 Din_27 n4825 VDD GND XOR2_X1
xU6795 n4838 n4839 n4833 VDD GND XOR2_X1
xU6796 n352 n4840 n4839 VDD GND XOR2_X1
xU6797 n4841 n4842 n4834 VDD GND XOR2_X1
xU6798 n4843 n4844 n4842 VDD GND XOR2_X1
xU6799 n4822 n4746 n4844 VDD GND XOR2_X1
xU6800 n4845 n375 n4746 VDD GND XOR2_X1
xU6801 n640 n381 n4843 VDD GND XOR2_X1
xU6802 n4846 n4847 n4841 VDD GND XOR2_X1
xU6803 n4848 n320 n4847 VDD GND XOR2_X1
xU6804 n4849 n4850 n4846 VDD GND XOR2_X1
xU6805 n707 Din_26 n4853 VDD GND XOR2_X1
xU6806 n4866 n4867 n4862 VDD GND XOR2_X1
xU6807 n4868 n4869 n4867 VDD GND XOR2_X1
xU6808 n379 n4870 n4869 VDD GND XOR2_X1
xU6809 n4871 n4872 n4866 VDD GND XOR2_X1
xU6810 n4873 n4816 n4872 VDD GND XOR2_X1
xU6811 n4874 n4875 n4816 VDD GND XOR2_X1
xU6812 n706 Din_25 n4878 VDD GND XOR2_X1
xU6813 n4891 n4892 n4887 VDD GND XOR2_X1
xU6814 n4893 n4894 n4892 VDD GND XOR2_X1
xU6815 n4895 n496 n4891 VDD GND XOR2_X1
xU6816 n705 Din_24 n4898 VDD GND XOR2_X1
xU6817 n4911 n4720 n4906 VDD GND XOR2_X1
xU6818 n4912 n4913 n4907 VDD GND XOR2_X1
xU6819 n4914 n4915 n4913 VDD GND XOR2_X1
xU6820 n4916 n4917 n4915 VDD GND XOR2_X1
xU6821 n4918 n4919 n4912 VDD GND XOR2_X1
xU6822 n4725 n4712 n4919 VDD GND XOR2_X1
xU6823 n704 Din_23 n4922 VDD GND XOR2_X1
xU6824 n4935 n4936 n4931 VDD GND XOR2_X1
xU6825 n4937 n4938 n4936 VDD GND XOR2_X1
xU6826 n631 n4914 n4938 VDD GND XOR2_X1
xU6827 n4939 n503 n4914 VDD GND XOR2_X1
xU6828 n4940 n4941 n4935 VDD GND XOR2_X1
xU6829 n4942 n382 n4940 VDD GND XOR2_X1
xU6830 n703 Din_22 n4945 VDD GND XOR2_X1
xU6831 n4958 n4959 n4953 VDD GND XOR2_X1
xU6832 n4960 n4961 n4959 VDD GND XOR2_X1
xU6833 n323 n4962 n4961 VDD GND XOR2_X1
xU6834 n636 n4963 n4958 VDD GND XOR2_X1
xU6835 n4964 n4965 n4963 VDD GND XOR2_X1
xU6836 n702 Din_21 n4968 VDD GND XOR2_X1
xU6837 n4981 n4982 n4977 VDD GND XOR2_X1
xU6838 n4983 n4984 n4982 VDD GND XOR2_X1
xU6839 n4985 n4986 n4984 VDD GND XOR2_X1
xU6840 n4987 n4988 n4983 VDD GND XOR2_X1
xU6841 n4989 n4990 n4981 VDD GND XOR2_X1
xU6842 n4991 n4795 n4990 VDD GND XOR2_X1
xU6843 n335 n4962 n4989 VDD GND XOR2_X1
xU6844 n701 Din_20 n4994 VDD GND XOR2_X1
xU6845 n5006 n5007 n5002 VDD GND XOR2_X1
xU6846 n5008 n5009 n5007 VDD GND XOR2_X1
xU6847 n5010 n5011 n5009 VDD GND XOR2_X1
xU6848 n5012 n4819 n5006 VDD GND XOR2_X1
xU6849 n5013 n4848 n4819 VDD GND XOR2_X1
xU6850 n4845 n5014 n5012 VDD GND XOR2_X1
xU6851 n700 Din_19 n5017 VDD GND XOR2_X1
xU6852 n640 n5030 n5025 VDD GND XOR2_X1
xU6853 n5031 n5032 n5026 VDD GND XOR2_X1
xU6854 n5033 n5034 n5032 VDD GND XOR2_X1
xU6855 n4916 n5035 n5034 VDD GND XOR2_X1
xU6856 n5014 n5036 n4916 VDD GND XOR2_X1
xU6857 n5037 n5038 n5031 VDD GND XOR2_X1
xU6858 n4942 n4850 n5038 VDD GND XOR2_X1
xU6859 n507 n4711 n5037 VDD GND XOR2_X1
xU6860 n699 Din_18 n5041 VDD GND XOR2_X1
xU6861 n5053 n5054 n5049 VDD GND XOR2_X1
xU6862 n5055 n5056 n5054 VDD GND XOR2_X1
xU6863 n5057 n320 n5056 VDD GND XOR2_X1
xU6864 n5010 n5058 n5053 VDD GND XOR2_X1
xU6865 n4893 n4986 n5058 VDD GND XOR2_X1
xU6866 n5059 n5060 n4893 VDD GND XOR2_X1
xU6867 n5061 n4988 n5060 VDD GND XOR2_X1
xU6868 n637 n4875 n4988 VDD GND XOR2_X1
xU6869 n5062 n5063 n5059 VDD GND XOR2_X1
xU6870 n4717 n4770 n5063 VDD GND XOR2_X1
xU6871 n5064 n498 n5010 VDD GND XOR2_X1
xU6872 n698 Din_17 n5067 VDD GND XOR2_X1
xU6873 n5080 n5081 n5076 VDD GND XOR2_X1
xU6874 n4911 n5082 n5081 VDD GND XOR2_X1
xU6875 n371 n342 n5082 VDD GND XOR2_X1
xU6876 n5083 n5084 n5080 VDD GND XOR2_X1
xU6877 n4986 n5085 n5084 VDD GND XOR2_X1
xU6878 n640 n5086 n4986 VDD GND XOR2_X1
xU6879 n697 Din_16 n5089 VDD GND XOR2_X1
xU6880 n5102 n5103 n5098 VDD GND XOR2_X1
xU6881 n4911 n5104 n5103 VDD GND XOR2_X1
xU6882 n4750 n4894 n5104 VDD GND XOR2_X1
xU6883 n356 n4712 n4894 VDD GND XOR2_X1
xU6884 n4792 n5105 n4712 VDD GND XOR2_X1
xU6885 n5106 n5107 n5102 VDD GND XOR2_X1
xU6886 n5108 n5109 n5107 VDD GND XOR2_X1
xU6887 n696 Din_15 n5112 VDD GND XOR2_X1
xU6888 n506 n4750 n5120 VDD GND XOR2_X1
xU6889 n5125 n5126 n5121 VDD GND XOR2_X1
xU6890 n4937 n5127 n5126 VDD GND XOR2_X1
xU6891 n5128 n5129 n5127 VDD GND XOR2_X1
xU6892 n4719 n5130 n4937 VDD GND XOR2_X1
xU6893 n4930 n5106 n5125 VDD GND XOR2_X1
xU6894 n5131 n5132 n5106 VDD GND XOR2_X1
xU6895 n4820 n5133 n4930 VDD GND XOR2_X1
xU6896 n695 Din_14 n5136 VDD GND XOR2_X1
xU6897 n5148 n5149 n5144 VDD GND XOR2_X1
xU6898 n5150 n5151 n5149 VDD GND XOR2_X1
xU6899 n4745 n380 n5151 VDD GND XOR2_X1
xU6900 n4792 n5152 n4745 VDD GND XOR2_X1
xU6901 n631 n5153 n5148 VDD GND XOR2_X1
xU6902 n504 n5013 n5153 VDD GND XOR2_X1
xU6903 n694 Din_13 n5156 VDD GND XOR2_X1
xU6904 n5169 n5170 n5165 VDD GND XOR2_X1
xU6905 n5171 n5172 n5170 VDD GND XOR2_X1
xU6906 n636 n5173 n5172 VDD GND XOR2_X1
xU6907 n5174 n5175 n5169 VDD GND XOR2_X1
xU6908 n335 n5176 n5175 VDD GND XOR2_X1
xU6909 n5177 n5178 n4771 VDD GND XOR2_X1
xU6910 n5179 n5180 n5178 VDD GND XOR2_X1
xU6911 n5181 n5182 n5177 VDD GND XOR2_X1
xU6912 n5183 n5184 n5181 VDD GND XOR2_X1
xU6913 n5185 n380 n5174 VDD GND XOR2_X1
xU6914 n693 Din_12 n5188 VDD GND XOR2_X1
xU6915 n5200 n5201 n5196 VDD GND XOR2_X1
xU6916 n5202 n5203 n5201 VDD GND XOR2_X1
xU6917 n5204 n5108 n5203 VDD GND XOR2_X1
xU6918 n4942 n5205 n5108 VDD GND XOR2_X1
xU6919 n5011 n5206 n5200 VDD GND XOR2_X1
xU6920 n4725 n5207 n5206 VDD GND XOR2_X1
xU6921 n4811 n507 n5011 VDD GND XOR2_X1
xU6922 n692 Din_11 n5210 VDD GND XOR2_X1
xU6923 n4942 n5223 n5218 VDD GND XOR2_X1
xU6924 n5224 n5225 n5219 VDD GND XOR2_X1
xU6925 n5035 n5226 n5225 VDD GND XOR2_X1
xU6926 n5227 n4871 n5226 VDD GND XOR2_X1
xU6927 n500 n356 n4871 VDD GND XOR2_X1
xU6928 n4840 n5229 n5035 VDD GND XOR2_X1
xU6929 n5230 n5231 n4840 VDD GND XOR2_X1
xU6930 n5109 n5030 n5224 VDD GND XOR2_X1
xU6931 n4718 n5232 n5030 VDD GND XOR2_X1
xU6932 n635 n4820 n4718 VDD GND XOR2_X1
xU6933 n691 Din_10 n5235 VDD GND XOR2_X1
xU6934 n5248 n5249 n5243 VDD GND XOR2_X1
xU6935 n5033 n5250 n5249 VDD GND XOR2_X1
xU6936 n4861 n5251 n5250 VDD GND XOR2_X1
xU6937 n4792 n4814 n4861 VDD GND XOR2_X1
xU6938 n5252 n5253 n4814 VDD GND XOR2_X1
xU6939 n5179 n5230 n4792 VDD GND XOR2_X1
xU6940 n5204 n5254 n5248 VDD GND XOR2_X1
xU6941 n5083 n5171 n5254 VDD GND XOR2_X1
xU6942 n381 n5085 n5171 VDD GND XOR2_X1
xU6943 n5255 n498 n5085 VDD GND XOR2_X1
xU6944 n5257 n5258 n5083 VDD GND XOR2_X1
xU6945 n5259 n5260 n5258 VDD GND XOR2_X1
xU6946 n4962 n4939 n5257 VDD GND XOR2_X1
xU6947 n5261 n5262 n5204 VDD GND XOR2_X1
xU6948 n690 Din_9 n5265 VDD GND XOR2_X1
xU6949 n5278 n5279 n5274 VDD GND XOR2_X1
xU6950 n5075 n5280 n5279 VDD GND XOR2_X1
xU6951 n4886 n4723 n5280 VDD GND XOR2_X1
xU6952 n381 n5281 n4723 VDD GND XOR2_X1
xU6953 n5086 n5282 n5036 VDD GND XOR2_X1
xU6954 n343 n5283 n4886 VDD GND XOR2_X1
xU6955 n5284 n5285 n5278 VDD GND XOR2_X1
xU6956 n689 Din_8 n5288 VDD GND XOR2_X1
xU6957 n5301 n5109 n5296 VDD GND XOR2_X1
xU6958 n5302 n5303 n5297 VDD GND XOR2_X1
xU6959 n5304 n5305 n5303 VDD GND XOR2_X1
xU6960 n5306 n5097 n5305 VDD GND XOR2_X1
xU6961 n5086 n5281 n5097 VDD GND XOR2_X1
xU6962 n5185 n5014 n5281 VDD GND XOR2_X1
xU6963 n5130 n5307 n5302 VDD GND XOR2_X1
xU6964 n382 n4911 n5307 VDD GND XOR2_X1
xU6965 n4985 n4822 n4911 VDD GND XOR2_X1
xU6966 n688 Din_7 n5310 VDD GND XOR2_X1
xU6967 n5205 n382 n5318 VDD GND XOR2_X1
xU6968 n5323 n5324 n5319 VDD GND XOR2_X1
xU6969 n5304 n5325 n5324 VDD GND XOR2_X1
xU6970 n4960 n4918 n5325 VDD GND XOR2_X1
xU6971 n4845 n5133 n4918 VDD GND XOR2_X1
xU6972 n5326 n5230 n5304 VDD GND XOR2_X1
xU6973 n4873 n5182 n5230 VDD GND XOR2_X1
xU6974 n5327 n5328 n5182 VDD GND XOR2_X1
xU6975 n5329 n5152 n5323 VDD GND XOR2_X1
xU6976 n5330 n5331 n5152 VDD GND XOR2_X1
xU6977 n352 n4750 n5329 VDD GND XOR2_X1
xU6978 n687 Din_6 n5334 VDD GND XOR2_X1
xU6979 n5301 n5129 n4960 VDD GND XOR2_X1
xU6980 n5346 n5176 n5129 VDD GND XOR2_X1
xU6981 n5347 n5348 n5176 VDD GND XOR2_X1
xU6982 n5349 n5350 n5342 VDD GND XOR2_X1
xU6983 n631 n5351 n5350 VDD GND XOR2_X1
xU6984 n377 n343 n5351 VDD GND XOR2_X1
xU6985 n5352 n5231 n4811 VDD GND XOR2_X1
xU6986 n5105 n5253 n5231 VDD GND XOR2_X1
xU6987 n4985 n4743 n4957 VDD GND XOR2_X1
xU6988 n5353 n4790 n4743 VDD GND XOR2_X1
xU6989 n5354 n5355 n4790 VDD GND XOR2_X1
xU6990 n5128 n5356 n5349 VDD GND XOR2_X1
xU6991 n4873 n5357 n5356 VDD GND XOR2_X1
xU6992 n5185 n4941 n5128 VDD GND XOR2_X1
xU6993 n5358 n4991 n4941 VDD GND XOR2_X1
xU6994 n5359 n5360 n4991 VDD GND XOR2_X1
xU6995 n686 Din_5 n5363 VDD GND XOR2_X1
xU6996 n5375 n5376 n4795 VDD GND XOR2_X1
xU6997 n5227 n5173 n5376 VDD GND XOR2_X1
xU6998 n5377 n5150 n5173 VDD GND XOR2_X1
xU6999 n5378 n5379 n5150 VDD GND XOR2_X1
xU7000 n5380 n5381 n5379 VDD GND XOR2_X1
xU7001 Dout_E_33 n5384 n5382 VDD GND XOR2_X1
xU7002 n5385 n5386 n5375 VDD GND XOR2_X1
xU7003 n5387 n5388 n5385 VDD GND XOR2_X1
xU7004 n5389 n5390 n5371 VDD GND XOR2_X1
xU7005 n5391 n5392 n5390 VDD GND XOR2_X1
xU7006 n4976 n5393 n5392 VDD GND XOR2_X1
xU7007 n5394 n5395 n4976 VDD GND XOR2_X1
xU7008 n4791 n4848 n5395 VDD GND XOR2_X1
xU7009 n639 n5396 n4791 VDD GND XOR2_X1
xU7010 n5398 n5399 n5397 VDD GND XOR2_X1
xU7011 n5400 n5401 n5399 VDD GND XOR2_X1
xU7012 Dout_E_113 n5404 n5402 VDD GND XOR2_X1
xU7013 n5405 n5406 n5394 VDD GND XOR2_X1
xU7014 n5407 n5408 n5405 VDD GND XOR2_X1
xU7015 n5164 n5409 n5389 VDD GND XOR2_X1
xU7016 n5331 n5180 n5409 VDD GND XOR2_X1
xU7017 n5357 n5410 n5180 VDD GND XOR2_X1
xU7018 n354 n5411 n5357 VDD GND XOR2_X1
xU7019 n5412 n5413 n5411 VDD GND XOR2_X1
xU7020 n363 n5416 n5414 VDD GND XOR2_X1
xU7021 n5418 n5419 n5331 VDD GND XOR2_X1
xU7022 n5420 n5421 n5164 VDD GND XOR2_X1
xU7023 n507 n4987 n5421 VDD GND XOR2_X1
xU7024 n4964 n5422 n4987 VDD GND XOR2_X1
xU7025 n5423 n5424 n4964 VDD GND XOR2_X1
xU7026 n5425 n5426 n5424 VDD GND XOR2_X1
xU7027 Dout_E_73 n5429 n5427 VDD GND XOR2_X1
xU7028 n5430 n5431 n5420 VDD GND XOR2_X1
xU7029 n5432 n5433 n5430 VDD GND XOR2_X1
xU7030 n685 Din_4 n5436 VDD GND XOR2_X1
xU7031 n5448 n5449 n5444 VDD GND XOR2_X1
xU7032 n5202 n5450 n5449 VDD GND XOR2_X1
xU7033 n5451 n5229 n5450 VDD GND XOR2_X1
xU7034 n5252 n5130 n5229 VDD GND XOR2_X1
xU7035 n352 n5205 n5130 VDD GND XOR2_X1
xU7036 n4768 n5227 n5202 VDD GND XOR2_X1
xU7037 n4817 n5452 n5448 VDD GND XOR2_X1
xU7038 n5105 n5352 n5452 VDD GND XOR2_X1
xU7039 n497 n5179 n4817 VDD GND XOR2_X1
xU7040 n684 Din_3 n5455 VDD GND XOR2_X1
xU7041 n5468 n4850 n5463 VDD GND XOR2_X1
xU7042 n5469 n5470 n4850 VDD GND XOR2_X1
xU7043 n5261 n5132 n5470 VDD GND XOR2_X1
xU7044 n375 n5282 n5468 VDD GND XOR2_X1
xU7045 n5471 n5472 n5205 VDD GND XOR2_X1
xU7046 n5473 n5380 n5472 VDD GND XOR2_X1
xU7047 n388 n5476 n5474 VDD GND XOR2_X1
xU7048 n5479 n5480 n5464 VDD GND XOR2_X1
xU7049 n5481 n5482 n5480 VDD GND XOR2_X1
xU7050 n5306 n5223 n5482 VDD GND XOR2_X1
xU7051 n5086 n4849 n5223 VDD GND XOR2_X1
xU7052 n5483 n5484 n4849 VDD GND XOR2_X1
xU7053 n5064 n503 n5484 VDD GND XOR2_X1
xU7054 n5228 n5105 n5306 VDD GND XOR2_X1
xU7055 n5330 n5410 n5105 VDD GND XOR2_X1
xU7056 n640 n4711 n5228 VDD GND XOR2_X1
xU7057 n379 n5232 n5481 VDD GND XOR2_X1
xU7058 n4874 n5494 n5232 VDD GND XOR2_X1
xU7059 n5495 n5496 n5479 VDD GND XOR2_X1
xU7060 n5179 n4845 n5496 VDD GND XOR2_X1
xU7061 n4820 n4942 n4845 VDD GND XOR2_X1
xU7062 n5425 n5497 n4942 VDD GND XOR2_X1
xU7063 n5498 n5499 n5497 VDD GND XOR2_X1
xU7064 Dout_E_73 n5504 n5502 VDD GND XOR2_X1
xU7065 n5400 n5505 n4820 VDD GND XOR2_X1
xU7066 n5506 n5507 n5505 VDD GND XOR2_X1
xU7067 n5512 n5513 n5510 VDD GND XOR2_X1
xU7068 n4719 n5326 n5179 VDD GND XOR2_X1
xU7069 n635 n352 n5495 VDD GND XOR2_X1
xU7070 n5412 n5514 n4821 VDD GND XOR2_X1
xU7071 n5515 n5516 n5514 VDD GND XOR2_X1
xU7072 n683 Din_2 n5523 VDD GND XOR2_X1
xU7073 n5301 n5451 n5057 VDD GND XOR2_X1
xU7074 n5261 n5535 n5451 VDD GND XOR2_X1
xU7075 n5537 n5538 n5531 VDD GND XOR2_X1
xU7076 n5393 n5539 n5538 VDD GND XOR2_X1
xU7077 n5033 n5285 n5539 VDD GND XOR2_X1
xU7078 n5540 n5541 n5285 VDD GND XOR2_X1
xU7079 n5542 n5543 n5541 VDD GND XOR2_X1
xU7080 n5544 n5131 n5540 VDD GND XOR2_X1
xU7081 n4985 n5008 n5033 VDD GND XOR2_X1
xU7082 n4874 n5545 n5008 VDD GND XOR2_X1
xU7083 n4749 n4848 n4985 VDD GND XOR2_X1
xU7084 n5133 n4717 n4848 VDD GND XOR2_X1
xU7085 n4770 n5406 n4749 VDD GND XOR2_X1
xU7086 n5062 n5548 n5406 VDD GND XOR2_X1
xU7087 Dout_E_113 n5553 n5551 VDD GND XOR2_X1
xU7088 n5282 n5284 n5393 VDD GND XOR2_X1
xU7089 n5535 n5262 n5284 VDD GND XOR2_X1
xU7090 n5554 n5555 n5537 VDD GND XOR2_X1
xU7091 n500 n5283 n5555 VDD GND XOR2_X1
xU7092 n5556 n5557 n5283 VDD GND XOR2_X1
xU7093 n4719 n5328 n5556 VDD GND XOR2_X1
xU7094 n5558 n5559 n5488 VDD GND XOR2_X1
xU7095 n367 n5562 n5560 VDD GND XOR2_X1
xU7096 n5185 n5207 n5247 VDD GND XOR2_X1
xU7097 n5064 n5255 n5207 VDD GND XOR2_X1
xU7098 n507 n5485 n5185 VDD GND XOR2_X1
xU7099 n4962 n5431 n5485 VDD GND XOR2_X1
xU7100 n5259 n5564 n5431 VDD GND XOR2_X1
xU7101 Dout_E_73 n5569 n5567 VDD GND XOR2_X1
xU7102 n4750 n4939 n5570 VDD GND XOR2_X1
xU7103 n5352 n4838 n5554 VDD GND XOR2_X1
xU7104 n4711 n5252 n4838 VDD GND XOR2_X1
xU7105 n682 Din_1 n5578 VDD GND XOR2_X1
xU7106 n5013 n5251 n4895 VDD GND XOR2_X1
xU7107 n5590 n5543 n5251 VDD GND XOR2_X1
xU7108 n5471 n5378 n5543 VDD GND XOR2_X1
xU7109 n5595 n5596 n5590 VDD GND XOR2_X1
xU7110 n5262 n5469 n5013 VDD GND XOR2_X1
xU7111 n4725 n5535 n5469 VDD GND XOR2_X1
xU7112 n5348 n5388 n5535 VDD GND XOR2_X1
xU7113 n5347 n5387 n5262 VDD GND XOR2_X1
xU7114 n5602 n5603 n5586 VDD GND XOR2_X1
xU7115 n5109 n5391 n5603 VDD GND XOR2_X1
xU7116 n4917 n4873 n5391 VDD GND XOR2_X1
xU7117 Dout_E_29 n5606 n5604 VDD GND XOR2_X1
xU7118 n378 n4711 n4917 VDD GND XOR2_X1
xU7119 n5608 n357 n5561 VDD GND XOR2_X1
xU7120 n5558 n5575 n5608 VDD GND XOR2_X1
xU7121 n5227 n5132 n5301 VDD GND XOR2_X1
xU7122 n380 n5386 n5132 VDD GND XOR2_X1
xU7123 n5542 n5596 n5386 VDD GND XOR2_X1
xU7124 n5475 n5597 n5600 VDD GND XOR2_X1
xU7125 n5614 n5615 n5597 VDD GND XOR2_X1
xU7126 Dout_E_33 n5592 n5613 VDD GND XOR2_X1
xU7127 n382 n5131 n5227 VDD GND XOR2_X1
xU7128 n4725 n5282 n5109 VDD GND XOR2_X1
xU7129 n5383 n5609 n5617 VDD GND XOR2_X1
xU7130 n5346 n5377 n4725 VDD GND XOR2_X1
xU7131 n5615 n5623 n5609 VDD GND XOR2_X1
xU7132 n5625 n5626 n5620 VDD GND XOR2_X1
xU7133 n5477 n5591 n5593 VDD GND XOR2_X1
xU7134 n5614 n5623 n5591 VDD GND XOR2_X1
xU7135 n5634 n5621 n5630 VDD GND XOR2_X1
xU7136 n5635 n5636 n5621 VDD GND XOR2_X1
xU7137 n5476 n5637 n5635 VDD GND XOR2_X1
xU7138 n5641 n5642 n5640 VDD GND XOR2_X1
xU7139 n5643 n5610 n5642 VDD GND XOR2_X1
xU7140 n5644 n5645 n5639 VDD GND XOR2_X1
xU7141 n5384 n5646 n5645 VDD GND XOR2_X1
xU7142 n5647 n5648 n5626 VDD GND XOR2_X1
xU7143 n5594 n5636 n5648 VDD GND XOR2_X1
xU7144 n5649 n5650 n5636 VDD GND XOR2_X1
xU7145 n5633 n5651 n5632 VDD GND XOR2_X1
xU7146 n5627 n5638 n5651 VDD GND XOR2_X1
xU7147 n5641 n5653 n5624 VDD GND XOR2_X1
xU7148 n5654 n5384 n5653 VDD GND XOR2_X1
xU7149 n5610 n5594 n5384 VDD GND XOR2_X1
xU7150 n5649 n5655 n5641 VDD GND XOR2_X1
xU7151 n386 n5476 n5656 VDD GND XOR2_X1
xU7152 n385 n5657 n5652 VDD GND XOR2_X1
xU7153 n5478 n5646 n5657 VDD GND XOR2_X1
xU7154 n5655 n5650 n5646 VDD GND XOR2_X1
xU7155 Dout_E_32 n5659 n5658 VDD GND XOR2_X1
xU7156 Dout_E_38 n5601 n5598 VDD GND XOR2_X1
xU7157 Dout_E_32 n5592 n5601 VDD GND XOR2_X1
xU7158 Dout_E_37 n5660 n5592 VDD GND XOR2_X1
xU7159 Dout_E_35 n391 n5661 VDD GND XOR2_X1
xU7160 Dout_E_33 n5662 n5536 VDD GND XOR2_X1
xU7161 Dout_E_37 Dout_E_39 n5478 VDD GND XOR2_X1
xU7162 n384 n5643 n5631 VDD GND XOR2_X1
xU7163 n5665 n5666 n5643 VDD GND XOR2_X1
xU7164 n5594 n5654 n5667 VDD GND XOR2_X1
xU7165 n5668 n5669 n5654 VDD GND XOR2_X1
xU7166 n5663 n5670 n5664 VDD GND XOR2_X1
xU7167 n5476 n5644 n5670 VDD GND XOR2_X1
xU7168 n387 n5665 n5644 VDD GND XOR2_X1
xU7169 Dout_E_36 n5672 n5671 VDD GND XOR2_X1
xU7170 n5674 n5660 n5476 VDD GND XOR2_X1
xU7171 n5669 n5675 n5663 VDD GND XOR2_X1
xU7172 n5659 n5677 n5676 VDD GND XOR2_X1
xU7173 Dout_E_39 Dout_E_34 n5677 VDD GND XOR2_X1
xU7174 n5662 n5659 n5599 VDD GND XOR2_X1
xU7175 n394 n388 n5659 VDD GND XOR2_X1
xU7176 n5678 n5679 n5633 VDD GND XOR2_X1
xU7177 n5674 n5647 n5679 VDD GND XOR2_X1
xU7178 n5673 n5666 n5647 VDD GND XOR2_X1
xU7179 Dout_E_35 n5681 n5629 VDD GND XOR2_X1
xU7180 Dout_E_34 n5681 n5680 VDD GND XOR2_X1
xU7181 n392 n395 n5681 VDD GND XOR2_X1
xU7182 n5610 n5672 n5616 VDD GND XOR2_X1
xU7183 Dout_E_33 n5660 n5672 VDD GND XOR2_X1
xU7184 Dout_E_39 n5594 n5660 VDD GND XOR2_X1
xU7185 Dout_E_34 Dout_E_35 n5594 VDD GND XOR2_X1
xU7186 Dout_E_37 n391 n5610 VDD GND XOR2_X1
xU7187 n392 Dout_E_38 n5674 VDD GND XOR2_X1
xU7188 Dout_E_39 n5637 n5678 VDD GND XOR2_X1
xU7189 n5668 n5675 n5637 VDD GND XOR2_X1
xU7190 Dout_E_33 n5684 n5622 VDD GND XOR2_X1
xU7191 Dout_E_32 n5686 n5685 VDD GND XOR2_X1
xU7192 Dout_E_38 Dout_E_35 n5686 VDD GND XOR2_X1
xU7193 n5662 n5684 n5618 VDD GND XOR2_X1
xU7194 n386 n392 n5684 VDD GND XOR2_X1
xU7195 Dout_E_34 Dout_E_37 n5662 VDD GND XOR2_X1
xU7196 n5075 n5687 n5602 VDD GND XOR2_X1
xU7197 n4870 n496 n5687 VDD GND XOR2_X1
xU7198 n4965 n5055 n5273 VDD GND XOR2_X1
xU7199 n5260 n5688 n5055 VDD GND XOR2_X1
xU7200 n4750 n5564 n5688 VDD GND XOR2_X1
xU7201 n5428 n5689 n5486 VDD GND XOR2_X1
xU7202 n5566 n514 n5429 VDD GND XOR2_X1
xU7203 n5498 n5423 n5260 VDD GND XOR2_X1
xU7204 n5256 n5483 n4965 VDD GND XOR2_X1
xU7205 n5014 n5255 n5483 VDD GND XOR2_X1
xU7206 n5360 n5432 n5255 VDD GND XOR2_X1
xU7207 n5358 n5422 n5014 VDD GND XOR2_X1
xU7208 n5695 n5696 n5689 VDD GND XOR2_X1
xU7209 n5500 n5571 n5692 VDD GND XOR2_X1
xU7210 n5696 n5698 n5571 VDD GND XOR2_X1
xU7211 n5359 n5433 n5256 VDD GND XOR2_X1
xU7212 n5704 n5705 n5699 VDD GND XOR2_X1
xU7213 n5706 n5707 n5705 VDD GND XOR2_X1
xU7214 n5503 n5568 n5565 VDD GND XOR2_X1
xU7215 n5695 n5698 n5568 VDD GND XOR2_X1
xU7216 n5713 n5714 n5704 VDD GND XOR2_X1
xU7217 n509 n5715 n5714 VDD GND XOR2_X1
xU7218 n5504 n5716 n5713 VDD GND XOR2_X1
xU7219 n5717 n5718 n5711 VDD GND XOR2_X1
xU7220 n5706 n5719 n5718 VDD GND XOR2_X1
xU7221 n512 n5721 n5710 VDD GND XOR2_X1
xU7222 n5715 n5722 n5721 VDD GND XOR2_X1
xU7223 n5723 n5724 n5720 VDD GND XOR2_X1
xU7224 n5725 n512 n5724 VDD GND XOR2_X1
xU7225 n514 n5727 n5723 VDD GND XOR2_X1
xU7226 n5729 n5730 n5717 VDD GND XOR2_X1
xU7227 n509 n5731 n5730 VDD GND XOR2_X1
xU7228 n510 n5732 n5709 VDD GND XOR2_X1
xU7229 n5719 n5707 n5732 VDD GND XOR2_X1
xU7230 n5726 n5734 n5712 VDD GND XOR2_X1
xU7231 n5729 n5735 n5734 VDD GND XOR2_X1
xU7232 n5715 n5728 n5729 VDD GND XOR2_X1
xU7233 Dout_E_72 n5504 n5736 VDD GND XOR2_X1
xU7234 n5737 n5566 n5726 VDD GND XOR2_X1
xU7235 n5738 n5739 n5733 VDD GND XOR2_X1
xU7236 n5740 n5501 n5739 VDD GND XOR2_X1
xU7237 n518 n520 n5501 VDD GND XOR2_X1
xU7238 n5727 n5737 n5738 VDD GND XOR2_X1
xU7239 Dout_E_75 n5742 n5741 VDD GND XOR2_X1
xU7240 Dout_E_73 n5743 n5563 VDD GND XOR2_X1
xU7241 Dout_E_72 n5745 n5744 VDD GND XOR2_X1
xU7242 Dout_E_78 n5708 n5693 VDD GND XOR2_X1
xU7243 Dout_E_72 n5569 n5708 VDD GND XOR2_X1
xU7244 Dout_E_77 n5746 n5569 VDD GND XOR2_X1
xU7245 n5748 n5722 n5700 VDD GND XOR2_X1
xU7246 n5749 n5750 n5722 VDD GND XOR2_X1
xU7247 n5728 n5735 n5748 VDD GND XOR2_X1
xU7248 n5751 n5752 n5735 VDD GND XOR2_X1
xU7249 n5753 n5725 n5747 VDD GND XOR2_X1
xU7250 n5754 n5749 n5725 VDD GND XOR2_X1
xU7251 Dout_E_76 n5756 n5755 VDD GND XOR2_X1
xU7252 n5504 n5740 n5753 VDD GND XOR2_X1
xU7253 n5751 n5757 n5740 VDD GND XOR2_X1
xU7254 n5745 n5759 n5758 VDD GND XOR2_X1
xU7255 Dout_E_79 Dout_E_74 n5759 VDD GND XOR2_X1
xU7256 n5743 n5745 n5701 VDD GND XOR2_X1
xU7257 n519 n513 n5745 VDD GND XOR2_X1
xU7258 n5742 n5746 n5504 VDD GND XOR2_X1
xU7259 n5760 n5761 n5703 VDD GND XOR2_X1
xU7260 n5716 n5731 n5761 VDD GND XOR2_X1
xU7261 n5754 n5750 n5731 VDD GND XOR2_X1
xU7262 Dout_E_75 n5763 n5697 VDD GND XOR2_X1
xU7263 Dout_E_74 n5763 n5762 VDD GND XOR2_X1
xU7264 n517 n520 n5763 VDD GND XOR2_X1
xU7265 n5566 n5756 n5572 VDD GND XOR2_X1
xU7266 Dout_E_73 n5746 n5756 VDD GND XOR2_X1
xU7267 n520 n5728 n5746 VDD GND XOR2_X1
xU7268 n515 Dout_E_75 n5728 VDD GND XOR2_X1
xU7269 Dout_E_77 n5742 n5566 VDD GND XOR2_X1
xU7270 n5752 n5757 n5716 VDD GND XOR2_X1
xU7271 Dout_E_73 n5766 n5694 VDD GND XOR2_X1
xU7272 n5743 n5766 n5487 VDD GND XOR2_X1
xU7273 n511 n517 n5766 VDD GND XOR2_X1
xU7274 Dout_E_74 Dout_E_77 n5743 VDD GND XOR2_X1
xU7275 Dout_E_72 n5768 n5767 VDD GND XOR2_X1
xU7276 Dout_E_78 Dout_E_75 n5768 VDD GND XOR2_X1
xU7277 n520 n5742 n5760 VDD GND XOR2_X1
xU7278 n517 n519 n5742 VDD GND XOR2_X1
xU7279 n5769 n5770 n4870 VDD GND XOR2_X1
xU7280 n4796 n5557 n5770 VDD GND XOR2_X1
xU7281 n5515 n5417 n5557 VDD GND XOR2_X1
xU7282 n5517 n5771 n5490 VDD GND XOR2_X1
xU7283 n5352 n5253 n4796 VDD GND XOR2_X1
xU7284 n5419 n5184 n5253 VDD GND XOR2_X1
xU7285 n355 n5559 n5605 VDD GND XOR2_X1
xU7286 n5418 n5183 n5352 VDD GND XOR2_X1
xU7287 n5327 n5326 n5769 VDD GND XOR2_X1
xU7288 n5776 n5558 n5771 VDD GND XOR2_X1
xU7289 n5784 n5785 n5779 VDD GND XOR2_X1
xU7290 n5786 n5787 n5785 VDD GND XOR2_X1
xU7291 n5789 n357 n5780 VDD GND XOR2_X1
xU7292 n5574 n5559 n5790 VDD GND XOR2_X1
xU7293 n5793 n5794 n5784 VDD GND XOR2_X1
xU7294 n5795 n5796 n5794 VDD GND XOR2_X1
xU7295 n5797 n5798 n5792 VDD GND XOR2_X1
xU7296 n5786 n5799 n5798 VDD GND XOR2_X1
xU7297 n5801 n5802 n5800 VDD GND XOR2_X1
xU7298 n5803 n5804 n5802 VDD GND XOR2_X1
xU7299 n362 n5562 n5801 VDD GND XOR2_X1
xU7300 n5776 n5774 n5789 VDD GND XOR2_X1
xU7301 n5806 n5807 n5797 VDD GND XOR2_X1
xU7302 n5808 n5795 n5807 VDD GND XOR2_X1
xU7303 n5809 n5810 n5795 VDD GND XOR2_X1
xU7304 Dout_E_25 n5773 n5806 VDD GND XOR2_X1
xU7305 n5812 n5813 n5811 VDD GND XOR2_X1
xU7306 n5814 n5815 n5813 VDD GND XOR2_X1
xU7307 n5778 n5816 n5805 VDD GND XOR2_X1
xU7308 n5787 n5799 n5816 VDD GND XOR2_X1
xU7309 n360 n5818 n5783 VDD GND XOR2_X1
xU7310 n5773 n5815 n5818 VDD GND XOR2_X1
xU7311 n5819 n5820 n5815 VDD GND XOR2_X1
xU7312 n5822 n5823 n5821 VDD GND XOR2_X1
xU7313 n5824 n5825 n5817 VDD GND XOR2_X1
xU7314 n5520 n5803 n5825 VDD GND XOR2_X1
xU7315 n5826 n5819 n5803 VDD GND XOR2_X1
xU7316 Dout_E_28 n5606 n5827 VDD GND XOR2_X1
xU7317 n5828 n5773 n5606 VDD GND XOR2_X1
xU7318 n5822 n5829 n5824 VDD GND XOR2_X1
xU7319 n5796 n5831 n5791 VDD GND XOR2_X1
xU7320 n5822 n5812 n5831 VDD GND XOR2_X1
xU7321 n5809 n5832 n5812 VDD GND XOR2_X1
xU7322 n363 n5834 n5833 VDD GND XOR2_X1
xU7323 Dout_E_31 Dout_E_24 n5834 VDD GND XOR2_X1
xU7324 Dout_E_24 n5772 n5781 VDD GND XOR2_X1
xU7325 n5823 n5562 n5796 VDD GND XOR2_X1
xU7326 n5793 n5835 n5830 VDD GND XOR2_X1
xU7327 n5822 n5804 n5835 VDD GND XOR2_X1
xU7328 n5810 n5832 n5804 VDD GND XOR2_X1
xU7329 n5836 n367 n5832 VDD GND XOR2_X1
xU7330 Dout_E_26 n5416 n5573 VDD GND XOR2_X1
xU7331 n365 n5814 n5837 VDD GND XOR2_X1
xU7332 Dout_E_25 n5839 n5838 VDD GND XOR2_X1
xU7333 n5839 n5772 n5775 VDD GND XOR2_X1
xU7334 n5518 n5773 n5772 VDD GND XOR2_X1
xU7335 Dout_E_31 Dout_E_29 n5518 VDD GND XOR2_X1
xU7336 n5828 n5841 n5840 VDD GND XOR2_X1
xU7337 n5841 n5416 n5777 VDD GND XOR2_X1
xU7338 n362 n367 n5416 VDD GND XOR2_X1
xU7339 Dout_E_26 Dout_E_30 n5841 VDD GND XOR2_X1
xU7340 n5829 Dout_E_31 n5793 VDD GND XOR2_X1
xU7341 n5842 n5843 n5778 VDD GND XOR2_X1
xU7342 n5828 n5808 n5843 VDD GND XOR2_X1
xU7343 n5826 n5820 n5808 VDD GND XOR2_X1
xU7344 Dout_E_26 n5845 n5844 VDD GND XOR2_X1
xU7345 Dout_E_27 n5845 n5491 VDD GND XOR2_X1
xU7346 n366 n369 n5845 VDD GND XOR2_X1
xU7347 n362 n5814 n5846 VDD GND XOR2_X1
xU7348 Dout_E_29 n5520 n5782 VDD GND XOR2_X1
xU7349 n5828 n363 n5520 VDD GND XOR2_X1
xU7350 n5814 n5773 n5562 VDD GND XOR2_X1
xU7351 Dout_E_26 Dout_E_27 n5773 VDD GND XOR2_X1
xU7352 Dout_E_31 Dout_E_25 n5828 VDD GND XOR2_X1
xU7353 n5814 n5847 n5842 VDD GND XOR2_X1
xU7354 n5829 n5823 n5847 VDD GND XOR2_X1
xU7355 n5849 n5850 n5607 VDD GND XOR2_X1
xU7356 n364 n367 n5849 VDD GND XOR2_X1
xU7357 Dout_E_27 n5839 n5848 VDD GND XOR2_X1
xU7358 n361 n368 n5839 VDD GND XOR2_X1
xU7359 n362 n5850 n5489 VDD GND XOR2_X1
xU7360 n361 n366 n5850 VDD GND XOR2_X1
xU7361 n367 n5814 n5788 VDD GND XOR2_X1
xU7362 n366 Dout_E_30 n5814 VDD GND XOR2_X1
xU7363 n4768 n4868 n5075 VDD GND XOR2_X1
xU7364 n5851 n5061 n4868 VDD GND XOR2_X1
xU7365 n5506 n5398 n5061 VDD GND XOR2_X1
xU7366 n5133 n5548 n5851 VDD GND XOR2_X1
xU7367 n5403 n5853 n5492 VDD GND XOR2_X1
xU7368 n4875 n5494 n4768 VDD GND XOR2_X1
xU7369 n4822 n637 n5494 VDD GND XOR2_X1
xU7370 n5355 n5408 n5545 VDD GND XOR2_X1
xU7371 n5353 n5396 n4822 VDD GND XOR2_X1
xU7372 n5858 n5859 n5853 VDD GND XOR2_X1
xU7373 n5508 n5547 n5852 VDD GND XOR2_X1
xU7374 n5858 n5861 n5547 VDD GND XOR2_X1
xU7375 n5354 n5407 n4875 VDD GND XOR2_X1
xU7376 n5867 n5868 n5862 VDD GND XOR2_X1
xU7377 n5869 n5870 n5868 VDD GND XOR2_X1
xU7378 n5511 n5552 n5549 VDD GND XOR2_X1
xU7379 n5861 n5859 n5552 VDD GND XOR2_X1
xU7380 n5876 n5877 n5867 VDD GND XOR2_X1
xU7381 n648 n5878 n5876 VDD GND XOR2_X1
xU7382 n5879 n5880 n5872 VDD GND XOR2_X1
xU7383 n5550 n5883 n5875 VDD GND XOR2_X1
xU7384 n646 n5884 n5883 VDD GND XOR2_X1
xU7385 n644 n5885 n5882 VDD GND XOR2_X1
xU7386 n5404 n641 n5885 VDD GND XOR2_X1
xU7387 n5887 n5888 n5880 VDD GND XOR2_X1
xU7388 n5889 n5877 n5888 VDD GND XOR2_X1
xU7389 n5890 n5891 n5877 VDD GND XOR2_X1
xU7390 n5866 n5892 n5874 VDD GND XOR2_X1
xU7391 n5881 n5870 n5892 VDD GND XOR2_X1
xU7392 n5404 n5894 n5873 VDD GND XOR2_X1
xU7393 n5895 n5884 n5894 VDD GND XOR2_X1
xU7394 n5896 n5890 n5884 VDD GND XOR2_X1
xU7395 n5513 n5898 n5897 VDD GND XOR2_X1
xU7396 n5899 Dout_E_112 n5898 VDD GND XOR2_X1
xU7397 n5550 n649 n5404 VDD GND XOR2_X1
xU7398 n642 n5900 n5893 VDD GND XOR2_X1
xU7399 n5509 n641 n5900 VDD GND XOR2_X1
xU7400 n5896 n5891 n5901 VDD GND XOR2_X1
xU7401 Dout_E_112 n5903 n5902 VDD GND XOR2_X1
xU7402 Dout_E_118 n5871 n5856 VDD GND XOR2_X1
xU7403 n5553 Dout_E_112 n5871 VDD GND XOR2_X1
xU7404 n648 Dout_E_117 n5553 VDD GND XOR2_X1
xU7405 Dout_E_115 n652 n5904 VDD GND XOR2_X1
xU7406 Dout_E_113 n5905 n5546 VDD GND XOR2_X1
xU7407 Dout_E_117 Dout_E_119 n5509 VDD GND XOR2_X1
xU7408 n5907 n5908 n5906 VDD GND XOR2_X1
xU7409 n5910 n646 n5863 VDD GND XOR2_X1
xU7410 n5912 n5913 n5911 VDD GND XOR2_X1
xU7411 n649 n5895 n5910 VDD GND XOR2_X1
xU7412 n5907 n5914 n5895 VDD GND XOR2_X1
xU7413 n5915 n5916 n5909 VDD GND XOR2_X1
xU7414 n5917 n5886 n5916 VDD GND XOR2_X1
xU7415 n5918 n5912 n5886 VDD GND XOR2_X1
xU7416 n653 n5512 n5919 VDD GND XOR2_X1
xU7417 n5907 n648 n5915 VDD GND XOR2_X1
xU7418 n5903 n5921 n5920 VDD GND XOR2_X1
xU7419 Dout_E_119 Dout_E_114 n5921 VDD GND XOR2_X1
xU7420 n5905 n5903 n5864 VDD GND XOR2_X1
xU7421 n655 n647 n5903 VDD GND XOR2_X1
xU7422 n5922 n5887 n5866 VDD GND XOR2_X1
xU7423 n5918 n5913 n5887 VDD GND XOR2_X1
xU7424 Dout_E_114 n5924 n5923 VDD GND XOR2_X1
xU7425 Dout_E_115 n5924 n5860 VDD GND XOR2_X1
xU7426 n653 n656 n5924 VDD GND XOR2_X1
xU7427 n5512 n5550 n5927 VDD GND XOR2_X1
xU7428 Dout_E_117 n652 n5550 VDD GND XOR2_X1
xU7429 n5899 Dout_E_113 n5512 VDD GND XOR2_X1
xU7430 n656 n649 n5899 VDD GND XOR2_X1
xU7431 n650 Dout_E_115 n5889 VDD GND XOR2_X1
xU7432 n656 n5878 n5922 VDD GND XOR2_X1
xU7433 n5914 n5917 n5878 VDD GND XOR2_X1
xU7434 n5908 n652 n5917 VDD GND XOR2_X1
xU7435 n653 Dout_E_118 n5513 VDD GND XOR2_X1
xU7436 Dout_E_113 n5928 n5857 VDD GND XOR2_X1
xU7437 n5905 n5928 n5493 VDD GND XOR2_X1
xU7438 n643 n653 n5928 VDD GND XOR2_X1
xU7439 Dout_E_114 Dout_E_117 n5905 VDD GND XOR2_X1
xU7440 Dout_E_112 n5930 n5929 VDD GND XOR2_X1
xU7441 Dout_E_118 Dout_E_115 n5930 VDD GND XOR2_X1
xU7442 n681 Din_0 n5934 VDD GND XOR2_X1
xU7443 \AES_Comp_ENCa/KrgX_63 n6166 n6390 VDD GND XOR2_X1
xU7444 n948 n5940 n6166 VDD GND XOR2_X1
xU7445 n6618 n6619 n5940 VDD GND XOR2_X1
xU7446 n6620 n6621 n6619 VDD GND XOR2_X1
xU7447 n6622 n6623 n6618 VDD GND XOR2_X1
xU7448 \AES_Comp_ENCa/KrgX_127 n6624 n6623 VDD GND XOR2_X1
xU7449 \AES_Comp_ENCa/KrgX_62 n6173 n6397 VDD GND XOR2_X1
xU7450 \AES_Comp_ENCa/KrgX_94 n5949 n6173 VDD GND XOR2_X1
xU7451 n6635 n6636 n5949 VDD GND XOR2_X1
xU7452 n6637 n6638 n6636 VDD GND XOR2_X1
xU7453 n6639 n979 n6635 VDD GND XOR2_X1
xU7454 \AES_Comp_ENCa/KrgX_61 n6180 n6404 VDD GND XOR2_X1
xU7455 \AES_Comp_ENCa/KrgX_93 n5956 n6180 VDD GND XOR2_X1
xU7456 n6651 n6652 n5956 VDD GND XOR2_X1
xU7457 n6620 n6653 n6652 VDD GND XOR2_X1
xU7458 n6654 n6655 n6653 VDD GND XOR2_X1
xU7459 n6658 n6659 n6651 VDD GND XOR2_X1
xU7460 n6660 \AES_Comp_ENCa/KrgX_125 n6658 VDD GND XOR2_X1
xU7461 \AES_Comp_ENCa/KrgX_60 n6187 n6411 VDD GND XOR2_X1
xU7462 n945 n5963 n6187 VDD GND XOR2_X1
xU7463 n6670 n6671 n5963 VDD GND XOR2_X1
xU7464 n6672 n6673 n6671 VDD GND XOR2_X1
xU7465 n6674 n6675 n6673 VDD GND XOR2_X1
xU7466 n6676 n6677 n6672 VDD GND XOR2_X1
xU7467 n6682 n6683 n6670 VDD GND XOR2_X1
xU7468 n6684 n6685 n6683 VDD GND XOR2_X1
xU7469 n857 n6688 n6686 VDD GND XOR2_X1
xU7470 n6689 \AES_Comp_ENCa/KrgX_124 n6682 VDD GND XOR2_X1
xU7471 \AES_Comp_ENCa/KrgX_59 n6194 n6418 VDD GND XOR2_X1
xU7472 \AES_Comp_ENCa/KrgX_91 n5970 n6194 VDD GND XOR2_X1
xU7473 n6699 n6700 n5970 VDD GND XOR2_X1
xU7474 n6701 n6702 n6700 VDD GND XOR2_X1
xU7475 n6705 n976 n6699 VDD GND XOR2_X1
xU7476 \AES_Comp_ENCa/KrgX_58 n6201 n6425 VDD GND XOR2_X1
xU7477 \AES_Comp_ENCa/KrgX_90 n5977 n6201 VDD GND XOR2_X1
xU7478 n6715 n6716 n5977 VDD GND XOR2_X1
xU7479 n6717 n6718 n6716 VDD GND XOR2_X1
xU7480 n6638 n6719 n6718 VDD GND XOR2_X1
xU7481 n6720 n6721 n6638 VDD GND XOR2_X1
xU7482 n6722 n6684 n6721 VDD GND XOR2_X1
xU7483 n857 n6725 n6723 VDD GND XOR2_X1
xU7484 n6728 n6729 n6717 VDD GND XOR2_X1
xU7485 n6732 n6733 n6715 VDD GND XOR2_X1
xU7486 n6734 n6735 n6733 VDD GND XOR2_X1
xU7487 n6622 n975 n6732 VDD GND XOR2_X1
xU7488 \AES_Comp_ENCa/KrgX_57 n6208 n6432 VDD GND XOR2_X1
xU7489 n942 n5984 n6208 VDD GND XOR2_X1
xU7490 n6747 n6748 n5984 VDD GND XOR2_X1
xU7491 n6620 n6749 n6748 VDD GND XOR2_X1
xU7492 n6734 n6675 n6620 VDD GND XOR2_X1
xU7493 n6729 n6750 n6675 VDD GND XOR2_X1
xU7494 n6751 n6637 n6750 VDD GND XOR2_X1
xU7495 n6754 n6755 n6729 VDD GND XOR2_X1
xU7496 \AES_Comp_ENCa/KrgX_17 n6759 n6757 VDD GND XOR2_X1
xU7497 n6760 n6761 n6747 VDD GND XOR2_X1
xU7498 n974 n6735 n6761 VDD GND XOR2_X1
xU7499 \AES_Comp_ENCa/KrgX_56 n6215 n6439 VDD GND XOR2_X1
xU7500 n941 n5991 n6215 VDD GND XOR2_X1
xU7501 n6778 n6779 n5991 VDD GND XOR2_X1
xU7502 n6702 n6780 n6779 VDD GND XOR2_X1
xU7503 n6781 n6674 n6780 VDD GND XOR2_X1
xU7504 n6782 n6705 n6674 VDD GND XOR2_X1
xU7505 n6785 n850 n6752 VDD GND XOR2_X1
xU7506 n6659 n6719 n6702 VDD GND XOR2_X1
xU7507 n849 n6621 n6719 VDD GND XOR2_X1
xU7508 n6660 n6689 n6621 VDD GND XOR2_X1
xU7509 n6654 n6676 n6749 VDD GND XOR2_X1
xU7510 n6724 n6758 n6756 VDD GND XOR2_X1
xU7511 n6785 n6796 n6758 VDD GND XOR2_X1
xU7512 n6797 n6798 n6778 VDD GND XOR2_X1
xU7513 n973 n6637 n6798 VDD GND XOR2_X1
xU7514 n851 n6799 n6736 VDD GND XOR2_X1
xU7515 n6764 n6796 n6800 VDD GND XOR2_X1
xU7516 n6720 n6755 n6797 VDD GND XOR2_X1
xU7517 n850 n6796 n6790 VDD GND XOR2_X1
xU7518 n6804 n6805 n6801 VDD GND XOR2_X1
xU7519 n848 n6799 n6792 VDD GND XOR2_X1
xU7520 n6808 n6763 n6799 VDD GND XOR2_X1
xU7521 n6802 n6812 n6810 VDD GND XOR2_X1
xU7522 n6807 n6813 n6812 VDD GND XOR2_X1
xU7523 n6816 n6817 n6814 VDD GND XOR2_X1
xU7524 n6818 n6819 n6816 VDD GND XOR2_X1
xU7525 n852 n6820 n6802 VDD GND XOR2_X1
xU7526 n6821 n6725 n6820 VDD GND XOR2_X1
xU7527 n6784 n6785 n6823 VDD GND XOR2_X1
xU7528 n6825 n6826 n6815 VDD GND XOR2_X1
xU7529 n6827 n6828 n6826 VDD GND XOR2_X1
xU7530 n6829 n6818 n6825 VDD GND XOR2_X1
xU7531 n853 n6830 n6805 VDD GND XOR2_X1
xU7532 n6831 n6828 n6830 VDD GND XOR2_X1
xU7533 n6832 n6833 n6828 VDD GND XOR2_X1
xU7534 n6834 n6835 n6817 VDD GND XOR2_X1
xU7535 n6809 n6836 n6824 VDD GND XOR2_X1
xU7536 n6806 n6813 n6836 VDD GND XOR2_X1
xU7537 n6819 n6838 n6803 VDD GND XOR2_X1
xU7538 n6839 n6822 n6838 VDD GND XOR2_X1
xU7539 n6832 n6840 n6822 VDD GND XOR2_X1
xU7540 n854 n6725 n6841 VDD GND XOR2_X1
xU7541 n6759 \AES_Comp_ENCa/KrgX_16 n6795 VDD GND XOR2_X1
xU7542 n6688 n6829 n6819 VDD GND XOR2_X1
xU7543 n6827 n859 n6688 VDD GND XOR2_X1
xU7544 n856 n6842 n6837 VDD GND XOR2_X1
xU7545 n6727 n6821 n6842 VDD GND XOR2_X1
xU7546 n6835 n6843 n6821 VDD GND XOR2_X1
xU7547 \AES_Comp_ENCa/KrgX_17 n6845 n6844 VDD GND XOR2_X1
xU7548 n6759 n6845 n6794 VDD GND XOR2_X1
xU7549 \AES_Comp_ENCa/KrgX_21 n6846 n6759 VDD GND XOR2_X1
xU7550 \AES_Comp_ENCa/KrgX_23 \AES_Comp_ENCa/KrgX_21 n6727 VDD GND XOR2_X1
xU7551 n6829 n6839 n6847 VDD GND XOR2_X1
xU7552 \AES_Comp_ENCa/KrgX_19 n863 n6848 VDD GND XOR2_X1
xU7553 \AES_Comp_ENCa/KrgX_21 n6849 n6762 VDD GND XOR2_X1
xU7554 n6851 n6852 n6811 VDD GND XOR2_X1
xU7555 n859 n6853 n6851 VDD GND XOR2_X1
xU7556 n6854 n6855 n6850 VDD GND XOR2_X1
xU7557 n6725 n6852 n6855 VDD GND XOR2_X1
xU7558 n6818 n6839 n6852 VDD GND XOR2_X1
xU7559 \AES_Comp_ENCa/KrgX_23 n6857 n6856 VDD GND XOR2_X1
xU7560 \AES_Comp_ENCa/KrgX_21 n6857 n6783 VDD GND XOR2_X1
xU7561 \AES_Comp_ENCa/KrgX_22 n6849 n6857 VDD GND XOR2_X1
xU7562 n860 n857 n6849 VDD GND XOR2_X1
xU7563 \AES_Comp_ENCa/KrgX_20 n6859 n6858 VDD GND XOR2_X1
xU7564 n6860 n6846 n6725 VDD GND XOR2_X1
xU7565 n6861 n6862 n6809 VDD GND XOR2_X1
xU7566 n6853 n6854 n6862 VDD GND XOR2_X1
xU7567 n855 n6843 n6854 VDD GND XOR2_X1
xU7568 \AES_Comp_ENCa/KrgX_17 n6863 n6791 VDD GND XOR2_X1
xU7569 n862 n6859 n6753 VDD GND XOR2_X1
xU7570 \AES_Comp_ENCa/KrgX_17 n6846 n6859 VDD GND XOR2_X1
xU7571 n867 n6831 n6846 VDD GND XOR2_X1
xU7572 n860 \AES_Comp_ENCa/KrgX_19 n6831 VDD GND XOR2_X1
xU7573 n865 n863 n6827 VDD GND XOR2_X1
xU7574 n6840 n6833 n6853 VDD GND XOR2_X1
xU7575 \AES_Comp_ENCa/KrgX_18 n6867 n6866 VDD GND XOR2_X1
xU7576 \AES_Comp_ENCa/KrgX_19 n6867 n6793 VDD GND XOR2_X1
xU7577 n864 n867 n6867 VDD GND XOR2_X1
xU7578 n6869 n6863 n6737 VDD GND XOR2_X1
xU7579 n854 n864 n6863 VDD GND XOR2_X1
xU7580 n860 n865 n6869 VDD GND XOR2_X1
xU7581 \AES_Comp_ENCa/KrgX_19 n6845 n6868 VDD GND XOR2_X1
xU7582 n854 n866 n6845 VDD GND XOR2_X1
xU7583 n867 n863 n6861 VDD GND XOR2_X1
xU7584 n864 \AES_Comp_ENCa/KrgX_22 n6860 VDD GND XOR2_X1
xU7585 \AES_Comp_ENCa/KrgX_55 n6222 n6446 VDD GND XOR2_X1
xU7586 \AES_Comp_ENCa/KrgX_87 n5998 n6222 VDD GND XOR2_X1
xU7587 n6879 n6880 n5998 VDD GND XOR2_X1
xU7588 n6881 n6882 n6880 VDD GND XOR2_X1
xU7589 n6883 n6884 n6879 VDD GND XOR2_X1
xU7590 n972 n6885 n6884 VDD GND XOR2_X1
xU7591 \AES_Comp_ENCa/KrgX_54 n6229 n6453 VDD GND XOR2_X1
xU7592 \AES_Comp_ENCa/KrgX_86 n6005 n6229 VDD GND XOR2_X1
xU7593 n6895 n6896 n6005 VDD GND XOR2_X1
xU7594 n6897 \AES_Comp_ENCa/KrgX_118 n6895 VDD GND XOR2_X1
xU7595 \AES_Comp_ENCa/KrgX_53 n6236 n6460 VDD GND XOR2_X1
xU7596 \AES_Comp_ENCa/KrgX_85 n6012 n6236 VDD GND XOR2_X1
xU7597 n6907 n6908 n6012 VDD GND XOR2_X1
xU7598 n6882 n6909 n6908 VDD GND XOR2_X1
xU7599 n6910 n970 n6907 VDD GND XOR2_X1
xU7600 \AES_Comp_ENCa/KrgX_52 n6243 n6467 VDD GND XOR2_X1
xU7601 \AES_Comp_ENCa/KrgX_84 n6019 n6243 VDD GND XOR2_X1
xU7602 n6920 n6921 n6019 VDD GND XOR2_X1
xU7603 n6922 n6923 n6921 VDD GND XOR2_X1
xU7604 n6924 n6925 n6923 VDD GND XOR2_X1
xU7605 n6926 n6927 n6920 VDD GND XOR2_X1
xU7606 n969 n6928 n6927 VDD GND XOR2_X1
xU7607 \AES_Comp_ENCa/KrgX_9 n6931 n6929 VDD GND XOR2_X1
xU7608 \AES_Comp_ENCa/KrgX_51 n6250 n6474 VDD GND XOR2_X1
xU7609 n936 n6026 n6250 VDD GND XOR2_X1
xU7610 n6941 n6942 n6026 VDD GND XOR2_X1
xU7611 n6943 \AES_Comp_ENCa/KrgX_115 n6941 VDD GND XOR2_X1
xU7612 \AES_Comp_ENCa/KrgX_50 n6257 n6481 VDD GND XOR2_X1
xU7613 n935 n6033 n6257 VDD GND XOR2_X1
xU7614 n6953 n6954 n6033 VDD GND XOR2_X1
xU7615 n6955 n6956 n6954 VDD GND XOR2_X1
xU7616 n6896 n6957 n6956 VDD GND XOR2_X1
xU7617 n6958 n6959 n6896 VDD GND XOR2_X1
xU7618 n6960 n6928 n6959 VDD GND XOR2_X1
xU7619 n840 n6963 n6961 VDD GND XOR2_X1
xU7620 n6966 n6967 n6955 VDD GND XOR2_X1
xU7621 n6968 n6969 n6953 VDD GND XOR2_X1
xU7622 n967 n6881 n6969 VDD GND XOR2_X1
xU7623 n6972 n6973 n6968 VDD GND XOR2_X1
xU7624 \AES_Comp_ENCa/KrgX_49 n6264 n6488 VDD GND XOR2_X1
xU7625 \AES_Comp_ENCa/KrgX_81 n6040 n6264 VDD GND XOR2_X1
xU7626 n6983 n6984 n6040 VDD GND XOR2_X1
xU7627 n6967 n6882 n6984 VDD GND XOR2_X1
xU7628 n6973 n6925 n6882 VDD GND XOR2_X1
xU7629 n8246 n6985 n6925 VDD GND XOR2_X1
xU7631 \AES_Comp_ENCa/KrgX_9 n6994 n6992 VDD GND XOR2_X1
xU7632 n6998 n6999 n6983 VDD GND XOR2_X1
xU7633 n7000 \AES_Comp_ENCa/KrgX_113 n6998 VDD GND XOR2_X1
xU7634 \AES_Comp_ENCa/KrgX_48 n6271 n6495 VDD GND XOR2_X1
xU7635 \AES_Comp_ENCa/KrgX_80 n6047 n6271 VDD GND XOR2_X1
xU7636 n7010 n7011 n6047 VDD GND XOR2_X1
xU7637 n6924 n6942 n7011 VDD GND XOR2_X1
xU7638 n6910 n6957 n6942 VDD GND XOR2_X1
xU7639 n6922 n6909 n6957 VDD GND XOR2_X1
xU7640 n6883 n7000 n6909 VDD GND XOR2_X1
xU7641 n836 n7013 n6993 VDD GND XOR2_X1
xU7642 n6885 n6999 n6922 VDD GND XOR2_X1
xU7643 n7021 n834 n6990 VDD GND XOR2_X1
xU7644 n7014 n7017 n7021 VDD GND XOR2_X1
xU7645 n7022 n6943 n6924 VDD GND XOR2_X1
xU7646 n7024 n6985 n7010 VDD GND XOR2_X1
xU7647 n6897 n6966 n6985 VDD GND XOR2_X1
xU7648 n835 n7013 n7018 VDD GND XOR2_X1
xU7649 n7026 n834 n6970 VDD GND XOR2_X1
xU7650 n6996 n7013 n7027 VDD GND XOR2_X1
xU7651 n7031 n7032 n7028 VDD GND XOR2_X1
xU7652 n7033 n7034 n7032 VDD GND XOR2_X1
xU7653 n7025 n6997 n7026 VDD GND XOR2_X1
xU7654 n6958 n965 n7024 VDD GND XOR2_X1
xU7655 n6964 n6989 n7015 VDD GND XOR2_X1
xU7656 n7014 n7025 n6989 VDD GND XOR2_X1
xU7657 n7030 n7041 n7036 VDD GND XOR2_X1
xU7658 n7033 n7042 n7041 VDD GND XOR2_X1
xU7659 n7044 n7045 n7039 VDD GND XOR2_X1
xU7660 n6991 n7046 n7045 VDD GND XOR2_X1
xU7661 n7047 n7048 n7044 VDD GND XOR2_X1
xU7662 n7049 n7050 n7043 VDD GND XOR2_X1
xU7663 n7048 n7051 n7049 VDD GND XOR2_X1
xU7664 n837 n7052 n7030 VDD GND XOR2_X1
xU7665 n7053 n6963 n7052 VDD GND XOR2_X1
xU7666 n7040 n7055 n7038 VDD GND XOR2_X1
xU7667 n7034 n7042 n7055 VDD GND XOR2_X1
xU7668 n7051 n7057 n7029 VDD GND XOR2_X1
xU7669 n7058 n7054 n7057 VDD GND XOR2_X1
xU7670 n7059 n7060 n7054 VDD GND XOR2_X1
xU7671 n6931 n7047 n7051 VDD GND XOR2_X1
xU7672 n6991 n7035 n6931 VDD GND XOR2_X1
xU7673 n7061 n7062 n7056 VDD GND XOR2_X1
xU7674 n6965 n7053 n7062 VDD GND XOR2_X1
xU7675 n7063 n7064 n7053 VDD GND XOR2_X1
xU7676 \AES_Comp_ENCa/KrgX_15 \AES_Comp_ENCa/KrgX_13 n6965 VDD GND XOR2_X1
xU7677 n7047 n7058 n7061 VDD GND XOR2_X1
xU7678 \AES_Comp_ENCa/KrgX_11 n843 n7065 VDD GND XOR2_X1
xU7679 \AES_Comp_ENCa/KrgX_13 n7066 n6995 VDD GND XOR2_X1
xU7680 n7068 n7069 n7037 VDD GND XOR2_X1
xU7681 n7035 n7070 n7068 VDD GND XOR2_X1
xU7682 n838 n7071 n7067 VDD GND XOR2_X1
xU7683 n7069 n6963 n7071 VDD GND XOR2_X1
xU7684 n7048 n7058 n7069 VDD GND XOR2_X1
xU7685 \AES_Comp_ENCa/KrgX_15 n7073 n7072 VDD GND XOR2_X1
xU7686 \AES_Comp_ENCa/KrgX_13 n7073 n7023 VDD GND XOR2_X1
xU7687 \AES_Comp_ENCa/KrgX_14 n7066 n7073 VDD GND XOR2_X1
xU7688 n841 n840 n7066 VDD GND XOR2_X1
xU7689 \AES_Comp_ENCa/KrgX_12 n7075 n7074 VDD GND XOR2_X1
xU7690 n7077 n7078 n7040 VDD GND XOR2_X1
xU7691 n7079 n7076 n7078 VDD GND XOR2_X1
xU7692 n7080 n7064 n7076 VDD GND XOR2_X1
xU7693 \AES_Comp_ENCa/KrgX_9 n7081 n7019 VDD GND XOR2_X1
xU7694 n847 n7070 n7077 VDD GND XOR2_X1
xU7695 n7060 n7082 n7070 VDD GND XOR2_X1
xU7696 \AES_Comp_ENCa/KrgX_11 n7084 n7083 VDD GND XOR2_X1
xU7697 n7085 n7081 n6971 VDD GND XOR2_X1
xU7698 n844 n839 n7081 VDD GND XOR2_X1
xU7699 n841 n845 n7085 VDD GND XOR2_X1
xU7700 n7050 n7086 n7031 VDD GND XOR2_X1
xU7701 n7035 n7046 n7086 VDD GND XOR2_X1
xU7702 n7059 n7082 n7046 VDD GND XOR2_X1
xU7703 \AES_Comp_ENCa/KrgX_11 n7088 n7016 VDD GND XOR2_X1
xU7704 \AES_Comp_ENCa/KrgX_10 n7088 n7087 VDD GND XOR2_X1
xU7705 n844 n847 n7088 VDD GND XOR2_X1
xU7706 n839 n6963 n7089 VDD GND XOR2_X1
xU7707 n7079 n7090 n6963 VDD GND XOR2_X1
xU7708 n6994 \AES_Comp_ENCa/KrgX_8 n7020 VDD GND XOR2_X1
xU7709 n7080 n7063 n7050 VDD GND XOR2_X1
xU7710 \AES_Comp_ENCa/KrgX_9 n7084 n7091 VDD GND XOR2_X1
xU7711 n6994 n7084 n7012 VDD GND XOR2_X1
xU7712 n846 n839 n7084 VDD GND XOR2_X1
xU7713 \AES_Comp_ENCa/KrgX_13 n7090 n6994 VDD GND XOR2_X1
xU7714 n6991 n7075 n6988 VDD GND XOR2_X1
xU7715 \AES_Comp_ENCa/KrgX_9 n7090 n7075 VDD GND XOR2_X1
xU7716 \AES_Comp_ENCa/KrgX_15 n7035 n7090 VDD GND XOR2_X1
xU7717 \AES_Comp_ENCa/KrgX_10 \AES_Comp_ENCa/KrgX_11 n7035 VDD GND XOR2_X1
xU7718 \AES_Comp_ENCa/KrgX_13 n843 n6991 VDD GND XOR2_X1
xU7719 n844 \AES_Comp_ENCa/KrgX_14 n7079 VDD GND XOR2_X1
xU7720 \AES_Comp_ENCa/KrgX_47 n6278 n6502 VDD GND XOR2_X1
xU7721 n932 n6054 n6278 VDD GND XOR2_X1
xU7722 n7103 n7104 n6054 VDD GND XOR2_X1
xU7723 n7105 n7106 n7104 VDD GND XOR2_X1
xU7724 n7107 n7108 n7103 VDD GND XOR2_X1
xU7725 n7109 \AES_Comp_ENCa/KrgX_111 n7107 VDD GND XOR2_X1
xU7726 \AES_Comp_ENCa/KrgX_46 n6285 n6509 VDD GND XOR2_X1
xU7727 \AES_Comp_ENCa/KrgX_78 n6061 n6285 VDD GND XOR2_X1
xU7728 n7119 n7120 n6061 VDD GND XOR2_X1
xU7729 n963 n7121 n7119 VDD GND XOR2_X1
xU7730 \AES_Comp_ENCa/KrgX_45 n6292 n6516 VDD GND XOR2_X1
xU7731 \AES_Comp_ENCa/KrgX_77 n6068 n6292 VDD GND XOR2_X1
xU7732 n7131 n7132 n6068 VDD GND XOR2_X1
xU7733 \AES_Comp_ENCa/KrgX_109 n7106 n7132 VDD GND XOR2_X1
xU7734 \AES_Comp_ENCa/KrgX_44 n6299 n6523 VDD GND XOR2_X1
xU7735 n929 n6075 n6299 VDD GND XOR2_X1
xU7736 n7142 n7143 n6075 VDD GND XOR2_X1
xU7737 n7144 n7145 n7143 VDD GND XOR2_X1
xU7738 n7146 n7147 n7142 VDD GND XOR2_X1
xU7739 n961 n7148 n7147 VDD GND XOR2_X1
xU7740 \AES_Comp_ENCa/KrgX_1 n7151 n7149 VDD GND XOR2_X1
xU7741 \AES_Comp_ENCa/KrgX_43 n6306 n6530 VDD GND XOR2_X1
xU7742 n928 n6082 n6306 VDD GND XOR2_X1
xU7743 n7161 n7162 n6082 VDD GND XOR2_X1
xU7744 \AES_Comp_ENCa/KrgX_107 n7131 n7162 VDD GND XOR2_X1
xU7745 \AES_Comp_ENCa/KrgX_42 n6313 n6537 VDD GND XOR2_X1
xU7746 \AES_Comp_ENCa/KrgX_74 n6089 n6313 VDD GND XOR2_X1
xU7747 n7172 n7173 n6089 VDD GND XOR2_X1
xU7748 n7174 n7175 n7173 VDD GND XOR2_X1
xU7749 n7176 n7177 n7175 VDD GND XOR2_X1
xU7750 n7178 n7179 n7177 VDD GND XOR2_X1
xU7751 n7121 n7180 n7176 VDD GND XOR2_X1
xU7752 n7148 n7181 n7121 VDD GND XOR2_X1
xU7753 n825 n7186 n7184 VDD GND XOR2_X1
xU7754 n7187 n7188 n7174 VDD GND XOR2_X1
xU7755 n959 n7108 n7188 VDD GND XOR2_X1
xU7756 n7191 n7192 n7187 VDD GND XOR2_X1
xU7757 \AES_Comp_ENCa/KrgX_41 n6320 n6544 VDD GND XOR2_X1
xU7758 n926 n6096 n6320 VDD GND XOR2_X1
xU7759 n7202 n7203 n6096 VDD GND XOR2_X1
xU7760 n7178 n7106 n7203 VDD GND XOR2_X1
xU7761 n7192 n7144 n7106 VDD GND XOR2_X1
xU7762 n7204 n7179 n7144 VDD GND XOR2_X1
xU7763 n7205 n7206 n7179 VDD GND XOR2_X1
xU7765 \AES_Comp_ENCa/KrgX_1 n7215 n7213 VDD GND XOR2_X1
xU7766 n7219 n7220 n7202 VDD GND XOR2_X1
xU7767 n958 n7221 n7220 VDD GND XOR2_X1
xU7768 \AES_Comp_ENCa/KrgX_40 n6327 n6551 VDD GND XOR2_X1
xU7769 \AES_Comp_ENCa/KrgX_72 n6103 n6327 VDD GND XOR2_X1
xU7770 n7231 n7232 n6103 VDD GND XOR2_X1
xU7771 n7131 n7145 n7232 VDD GND XOR2_X1
xU7772 n7233 n7161 n7145 VDD GND XOR2_X1
xU7773 n7234 n7180 n7161 VDD GND XOR2_X1
xU7774 n7105 n7219 n7180 VDD GND XOR2_X1
xU7775 n7239 n7240 n7211 VDD GND XOR2_X1
xU7776 n7241 n7172 n7131 VDD GND XOR2_X1
xU7777 n7109 n7221 n7172 VDD GND XOR2_X1
xU7778 n7243 n7240 n7214 VDD GND XOR2_X1
xU7779 n7247 n7248 n7207 VDD GND XOR2_X1
xU7780 n7249 n7120 n7231 VDD GND XOR2_X1
xU7781 n7212 n7191 n7120 VDD GND XOR2_X1
xU7782 n7247 n7251 n7244 VDD GND XOR2_X1
xU7783 n7240 n7235 n7247 VDD GND XOR2_X1
xU7784 n7255 n7256 n7252 VDD GND XOR2_X1
xU7785 n7257 n7258 n7256 VDD GND XOR2_X1
xU7786 n7251 n7248 n7189 VDD GND XOR2_X1
xU7787 n7243 n7217 n7248 VDD GND XOR2_X1
xU7788 n7239 n7218 n7251 VDD GND XOR2_X1
xU7789 n7262 n7263 n7255 VDD GND XOR2_X1
xU7790 n7264 n7265 n7263 VDD GND XOR2_X1
xU7791 n832 n7266 n7262 VDD GND XOR2_X1
xU7792 n7206 n957 n7249 VDD GND XOR2_X1
xU7793 n7239 n7243 n7236 VDD GND XOR2_X1
xU7794 n7267 n7253 n7259 VDD GND XOR2_X1
xU7795 n7268 n7269 n7253 VDD GND XOR2_X1
xU7796 n7250 n7270 n7269 VDD GND XOR2_X1
xU7797 n7271 n7258 n7267 VDD GND XOR2_X1
xU7798 n7265 n7273 n7272 VDD GND XOR2_X1
xU7799 n7274 n7186 n7273 VDD GND XOR2_X1
xU7800 n7275 n7276 n7265 VDD GND XOR2_X1
xU7801 n7274 n7278 n7277 VDD GND XOR2_X1
xU7802 n7266 n7250 n7278 VDD GND XOR2_X1
xU7803 n7279 n7280 n7266 VDD GND XOR2_X1
xU7804 n7281 n7282 n7274 VDD GND XOR2_X1
xU7805 n7260 n7283 n7261 VDD GND XOR2_X1
xU7806 n7257 n7271 n7283 VDD GND XOR2_X1
xU7807 n7270 n7285 n7254 VDD GND XOR2_X1
xU7808 n7286 n7208 n7285 VDD GND XOR2_X1
xU7809 n7287 n7280 n7270 VDD GND XOR2_X1
xU7810 \AES_Comp_ENCa/KrgX_3 n7289 n7245 VDD GND XOR2_X1
xU7811 \AES_Comp_ENCa/KrgX_2 n7289 n7288 VDD GND XOR2_X1
xU7812 n829 n832 n7289 VDD GND XOR2_X1
xU7813 n7151 n7290 n7284 VDD GND XOR2_X1
xU7814 n7286 n7268 n7290 VDD GND XOR2_X1
xU7815 n7275 n7291 n7268 VDD GND XOR2_X1
xU7816 n7208 n7294 n7210 VDD GND XOR2_X1
xU7817 n7281 n7295 n7286 VDD GND XOR2_X1
xU7818 \AES_Comp_ENCa/KrgX_4 n7294 n7296 VDD GND XOR2_X1
xU7819 \AES_Comp_ENCa/KrgX_1 n7297 n7294 VDD GND XOR2_X1
xU7820 n7300 n7301 n7299 VDD GND XOR2_X1
xU7821 n7302 n7151 n7301 VDD GND XOR2_X1
xU7822 n7208 n7250 n7151 VDD GND XOR2_X1
xU7823 \AES_Comp_ENCa/KrgX_5 n828 n7208 VDD GND XOR2_X1
xU7824 n7182 n7303 n7298 VDD GND XOR2_X1
xU7825 n7304 n7300 n7303 VDD GND XOR2_X1
xU7826 n7282 n7295 n7300 VDD GND XOR2_X1
xU7827 \AES_Comp_ENCa/KrgX_3 n828 n7305 VDD GND XOR2_X1
xU7828 \AES_Comp_ENCa/KrgX_1 n7306 n7216 VDD GND XOR2_X1
xU7829 n7308 n7309 n7307 VDD GND XOR2_X1
xU7830 \AES_Comp_ENCa/KrgX_7 \AES_Comp_ENCa/KrgX_2 n7309 VDD GND XOR2_X1
xU7831 n7308 n7306 n7238 VDD GND XOR2_X1
xU7832 \AES_Comp_ENCa/KrgX_6 \AES_Comp_ENCa/KrgX_1 n7308 VDD GND XOR2_X1
xU7833 n830 \AES_Comp_ENCa/KrgX_7 n7182 VDD GND XOR2_X1
xU7834 n822 n7310 n7260 VDD GND XOR2_X1
xU7835 n7186 n7302 n7310 VDD GND XOR2_X1
xU7836 n7287 n7279 n7302 VDD GND XOR2_X1
xU7837 n7312 n7306 n7190 VDD GND XOR2_X1
xU7838 n826 n830 n7306 VDD GND XOR2_X1
xU7839 \AES_Comp_ENCa/KrgX_3 n7313 n7311 VDD GND XOR2_X1
xU7840 n824 n7186 n7314 VDD GND XOR2_X1
xU7841 n7215 \AES_Comp_ENCa/KrgX_0 n7246 VDD GND XOR2_X1
xU7842 n7264 n7297 n7186 VDD GND XOR2_X1
xU7843 n829 \AES_Comp_ENCa/KrgX_6 n7264 VDD GND XOR2_X1
xU7844 n7291 n7276 n7304 VDD GND XOR2_X1
xU7845 \AES_Comp_ENCa/KrgX_1 n7312 n7237 VDD GND XOR2_X1
xU7846 \AES_Comp_ENCa/KrgX_0 \AES_Comp_ENCa/KrgX_4 n7312 VDD GND XOR2_X1
xU7847 \AES_Comp_ENCa/KrgX_1 n7313 n7315 VDD GND XOR2_X1
xU7848 n7215 n7313 n7242 VDD GND XOR2_X1
xU7849 n824 n831 n7313 VDD GND XOR2_X1
xU7850 \AES_Comp_ENCa/KrgX_5 n7297 n7215 VDD GND XOR2_X1
xU7851 \AES_Comp_ENCa/KrgX_7 n7250 n7297 VDD GND XOR2_X1
xU7852 \AES_Comp_ENCa/KrgX_2 \AES_Comp_ENCa/KrgX_3 n7250 VDD GND XOR2_X1
xU7853 \AES_Comp_ENCa/KrgX_39 n6334 n6558 VDD GND XOR2_X1
xU7854 n924 n6110 n6334 VDD GND XOR2_X1
xU7855 n7325 n7326 n6110 VDD GND XOR2_X1
xU7856 n7327 n7328 n7326 VDD GND XOR2_X1
xU7857 n7329 \AES_Comp_ENCa/KrgX_103 n7325 VDD GND XOR2_X1
xU7858 \AES_Comp_ENCa/KrgX_38 n6341 n6565 VDD GND XOR2_X1
xU7859 \AES_Comp_ENCa/KrgX_70 n6117 n6341 VDD GND XOR2_X1
xU7860 n7339 n7340 n6117 VDD GND XOR2_X1
xU7861 n7341 \AES_Comp_ENCa/KrgX_102 n7339 VDD GND XOR2_X1
xU7862 \AES_Comp_ENCa/KrgX_37 n6348 n6572 VDD GND XOR2_X1
xU7863 \AES_Comp_ENCa/KrgX_69 n6124 n6348 VDD GND XOR2_X1
xU7864 n7351 n7352 n6124 VDD GND XOR2_X1
xU7865 n7353 n7327 n7352 VDD GND XOR2_X1
xU7866 n7354 n7355 n7351 VDD GND XOR2_X1
xU7867 n7356 n954 n7354 VDD GND XOR2_X1
xU7868 \AES_Comp_ENCa/KrgX_36 n6355 n6579 VDD GND XOR2_X1
xU7869 n921 n6131 n6355 VDD GND XOR2_X1
xU7870 n7366 n7367 n6131 VDD GND XOR2_X1
xU7871 n7368 n7369 n7367 VDD GND XOR2_X1
xU7872 n7370 n7371 n7369 VDD GND XOR2_X1
xU7873 n7373 n876 n7372 VDD GND XOR2_X1
xU7874 n7375 n7376 n7366 VDD GND XOR2_X1
xU7875 n7377 n7378 n7376 VDD GND XOR2_X1
xU7876 n7379 \AES_Comp_ENCa/KrgX_100 n7375 VDD GND XOR2_X1
xU7877 \AES_Comp_ENCa/KrgX_35 n6362 n6586 VDD GND XOR2_X1
xU7878 n920 n6138 n6362 VDD GND XOR2_X1
xU7879 n7389 n7390 n6138 VDD GND XOR2_X1
xU7880 n7391 \AES_Comp_ENCa/KrgX_99 n7389 VDD GND XOR2_X1
xU7881 \AES_Comp_ENCa/KrgX_34 n6369 n6593 VDD GND XOR2_X1
xU7882 n919 n6145 n6369 VDD GND XOR2_X1
xU7883 n7401 n7402 n6145 VDD GND XOR2_X1
xU7884 n7403 n7404 n7402 VDD GND XOR2_X1
xU7885 n7340 n7405 n7404 VDD GND XOR2_X1
xU7886 n7406 n7407 n7340 VDD GND XOR2_X1
xU7887 n7408 n7377 n7407 VDD GND XOR2_X1
xU7888 n876 n7411 n7409 VDD GND XOR2_X1
xU7889 n7414 n7415 n7403 VDD GND XOR2_X1
xU7890 n7416 n7417 n7401 VDD GND XOR2_X1
xU7891 n951 n7329 n7417 VDD GND XOR2_X1
xU7892 n7420 n7421 n7416 VDD GND XOR2_X1
xU7893 \AES_Comp_ENCa/KrgX_33 n6376 n6600 VDD GND XOR2_X1
xU7894 \AES_Comp_ENCa/KrgX_65 n6152 n6376 VDD GND XOR2_X1
xU7895 n7431 n7432 n6152 VDD GND XOR2_X1
xU7896 n7327 n7433 n7432 VDD GND XOR2_X1
xU7897 n7421 n7371 n7327 VDD GND XOR2_X1
xU7898 n8248 n7434 n7371 VDD GND XOR2_X1
xU7900 \AES_Comp_ENCa/KrgX_25 n7441 n7440 VDD GND XOR2_X1
xU7901 n7415 n950 n7431 VDD GND XOR2_X1
xU7902 \AES_Comp_ENCa/KrgX_32 n6383 n6607 VDD GND XOR2_X1
xU7903 \AES_Comp_ENCa/KrgX_64 n6159 n6383 VDD GND XOR2_X1
xU7904 n7457 n7458 n6159 VDD GND XOR2_X1
xU7905 n7368 n7390 n7458 VDD GND XOR2_X1
xU7906 n7355 n7405 n7390 VDD GND XOR2_X1
xU7907 n869 n7328 n7405 VDD GND XOR2_X1
xU7908 n7356 n7379 n7328 VDD GND XOR2_X1
xU7909 n7353 n7378 n7433 VDD GND XOR2_X1
xU7910 n7410 n871 n7439 VDD GND XOR2_X1
xU7911 n7466 n7467 n7465 VDD GND XOR2_X1
xU7912 n7470 n7391 n7368 VDD GND XOR2_X1
xU7913 n7472 n7434 n7457 VDD GND XOR2_X1
xU7914 n7341 n7414 n7434 VDD GND XOR2_X1
xU7915 n7374 n7459 n7418 VDD GND XOR2_X1
xU7916 n7466 n7473 n7459 VDD GND XOR2_X1
xU7917 n7477 n7478 n7474 VDD GND XOR2_X1
xU7918 n7479 n7480 n7478 VDD GND XOR2_X1
xU7919 n7406 n949 n7472 VDD GND XOR2_X1
xU7920 n7412 n870 n7461 VDD GND XOR2_X1
xU7921 n7473 n7467 n7438 VDD GND XOR2_X1
xU7922 n7476 n7486 n7483 VDD GND XOR2_X1
xU7923 n7479 n7487 n7486 VDD GND XOR2_X1
xU7924 n7489 n7490 n7482 VDD GND XOR2_X1
xU7925 n7491 n7492 n7490 VDD GND XOR2_X1
xU7926 n7493 n7494 n7489 VDD GND XOR2_X1
xU7927 n7495 n7496 n7488 VDD GND XOR2_X1
xU7928 n7494 n7497 n7496 VDD GND XOR2_X1
xU7929 n7498 n7499 n7476 VDD GND XOR2_X1
xU7930 n7500 n7411 n7499 VDD GND XOR2_X1
xU7931 n7497 n7501 n7477 VDD GND XOR2_X1
xU7932 n7502 n7491 n7501 VDD GND XOR2_X1
xU7933 n7503 n7504 n7491 VDD GND XOR2_X1
xU7934 n7505 n7506 n7497 VDD GND XOR2_X1
xU7935 n7485 n7507 n7481 VDD GND XOR2_X1
xU7936 n7480 n7487 n7507 VDD GND XOR2_X1
xU7937 n7495 n7510 n7509 VDD GND XOR2_X1
xU7938 n7511 n7498 n7510 VDD GND XOR2_X1
xU7939 n7503 n7512 n7498 VDD GND XOR2_X1
xU7940 n875 n7411 n7513 VDD GND XOR2_X1
xU7941 n7441 \AES_Comp_ENCa/KrgX_24 n7464 VDD GND XOR2_X1
xU7942 n7373 n7493 n7495 VDD GND XOR2_X1
xU7943 n881 n877 n7373 VDD GND XOR2_X1
xU7944 n7514 n7515 n7508 VDD GND XOR2_X1
xU7945 n7413 n7500 n7515 VDD GND XOR2_X1
xU7946 n7506 n7516 n7500 VDD GND XOR2_X1
xU7947 \AES_Comp_ENCa/KrgX_25 n7518 n7517 VDD GND XOR2_X1
xU7948 n7441 n7518 n7463 VDD GND XOR2_X1
xU7949 \AES_Comp_ENCa/KrgX_29 n7519 n7441 VDD GND XOR2_X1
xU7950 \AES_Comp_ENCa/KrgX_31 \AES_Comp_ENCa/KrgX_29 n7413 VDD GND XOR2_X1
xU7951 n7493 n7511 n7514 VDD GND XOR2_X1
xU7952 n879 n7521 n7520 VDD GND XOR2_X1
xU7953 \AES_Comp_ENCa/KrgX_29 n7522 n7442 VDD GND XOR2_X1
xU7954 n7523 n7524 n7484 VDD GND XOR2_X1
xU7955 n877 n7525 n7524 VDD GND XOR2_X1
xU7956 n7527 n7528 n7526 VDD GND XOR2_X1
xU7957 n7411 n7525 n7528 VDD GND XOR2_X1
xU7958 n7494 n7511 n7525 VDD GND XOR2_X1
xU7959 \AES_Comp_ENCa/KrgX_31 n7530 n7529 VDD GND XOR2_X1
xU7960 \AES_Comp_ENCa/KrgX_29 n7530 n7471 VDD GND XOR2_X1
xU7961 \AES_Comp_ENCa/KrgX_30 n7522 n7530 VDD GND XOR2_X1
xU7962 n878 n876 n7522 VDD GND XOR2_X1
xU7963 \AES_Comp_ENCa/KrgX_28 n7532 n7531 VDD GND XOR2_X1
xU7964 n7521 n7519 n7411 VDD GND XOR2_X1
xU7965 n7533 n7534 n7485 VDD GND XOR2_X1
xU7966 n7527 n7523 n7534 VDD GND XOR2_X1
xU7967 n7512 n7504 n7523 VDD GND XOR2_X1
xU7968 \AES_Comp_ENCa/KrgX_26 n7536 n7535 VDD GND XOR2_X1
xU7969 \AES_Comp_ENCa/KrgX_27 n7536 n7462 VDD GND XOR2_X1
xU7970 n880 n884 n7536 VDD GND XOR2_X1
xU7971 n7538 n7539 n7419 VDD GND XOR2_X1
xU7972 n878 n882 n7538 VDD GND XOR2_X1
xU7973 \AES_Comp_ENCa/KrgX_27 n7518 n7537 VDD GND XOR2_X1
xU7974 n875 n883 n7518 VDD GND XOR2_X1
xU7975 n7505 n7516 n7527 VDD GND XOR2_X1
xU7976 \AES_Comp_ENCa/KrgX_25 n7539 n7460 VDD GND XOR2_X1
xU7977 n875 n880 n7539 VDD GND XOR2_X1
xU7978 n7492 n7532 n7437 VDD GND XOR2_X1
xU7979 \AES_Comp_ENCa/KrgX_25 n7519 n7532 VDD GND XOR2_X1
xU7980 n884 n7502 n7519 VDD GND XOR2_X1
xU7981 n878 \AES_Comp_ENCa/KrgX_27 n7502 VDD GND XOR2_X1
xU7982 \AES_Comp_ENCa/KrgX_29 n7521 n7492 VDD GND XOR2_X1
xU7983 n884 n7521 n7533 VDD GND XOR2_X1
xU7984 \AES_Comp_ENCa/KrgX_28 n883 n7521 VDD GND XOR2_X1
xAES_Comp_ENCa/KrgX_reg_1 n8100 CLK \AES_Comp_ENCa/KrgX_1 n825 VDD GND DFF_X1
xU7985 n136 n7573 n8245 VDD GND AND2_X1
xU7986 n4375 n613 VDD GND INV_X1
xU7987 n4242 n282 VDD GND INV_X1
xU7988 n5025 n634 VDD GND INV_X1
xU7989 n5219 n330 VDD GND INV_X1
xU7990 n1583 n172 VDD GND INV_X1
xU7991 n5296 n370 VDD GND INV_X1
xU7992 n1381 n400 VDD GND INV_X1
xU7993 n2325 n548 VDD GND INV_X1
xU7994 n2283 n421 VDD GND INV_X1
xU7995 n1480 n397 VDD GND INV_X1
xU7996 n1146 n660 VDD GND INV_X1
xU7997 n3776 n478 VDD GND INV_X1
xU7998 n1240 n523 VDD GND INV_X1
xU7999 n4957 n631 VDD GND INV_X1
xU8000 n2738 n203 VDD GND INV_X1
xU8001 n1040 n661 VDD GND INV_X1
xU8002 n3570 n450 VDD GND INV_X1
xU8003 n3763 n262 VDD GND INV_X1
xU8004 n4960 n374 VDD GND INV_X1
xU8005 n4745 n323 VDD GND INV_X1
xU8006 n3528 n603 VDD GND INV_X1
xU8007 n3504 n447 VDD GND INV_X1
xU8008 n1089 n664 VDD GND INV_X1
xU8009 n3701 n269 VDD GND INV_X1
xU8010 n5013 n372 VDD GND INV_X1
xU8011 n4965 n497 VDD GND INV_X1
xU8012 n2482 n424 VDD GND INV_X1
xU8013 n4861 n320 VDD GND INV_X1
xU8014 n1734 n179 VDD GND INV_X1
xU8015 n5128 n499 VDD GND INV_X1
xU8016 n2258 n549 VDD GND INV_X1
xU8017 n3728 n602 VDD GND INV_X1
xU8018 n5033 n632 VDD GND INV_X1
xU8019 n4811 n343 VDD GND INV_X1
xU8020 n4768 n630 VDD GND INV_X1
xU8021 n5057 n379 VDD GND INV_X1
xU8022 n1428 n398 VDD GND INV_X1
xU8023 n1283 n522 VDD GND INV_X1
xU8024 n4098 n471 VDD GND INV_X1
xU8025 n1612 n161 VDD GND INV_X1
xU8026 n5247 n500 VDD GND INV_X1
xU8027 n2384 n550 VDD GND INV_X1
xU8028 n5301 n378 VDD GND INV_X1
xU8029 n2580 n426 VDD GND INV_X1
xU8030 n1335 n524 VDD GND INV_X1
xU8031 n4025 n454 VDD GND INV_X1
xU8032 n2978 n580 VDD GND INV_X1
xU8033 n1196 n153 VDD GND INV_X1
xU8034 n2224 n551 VDD GND INV_X1
xU8035 n2912 n582 VDD GND INV_X1
xU8036 n2634 n209 VDD GND INV_X1
xU8037 n3670 n281 VDD GND INV_X1
xU8038 n1191 n525 VDD GND INV_X1
xU8039 n5097 n501 VDD GND INV_X1
xU8040 n5036 n381 VDD GND INV_X1
xU8041 n3693 n296 VDD GND INV_X1
xU8042 n4227 n473 VDD GND INV_X1
xU8043 n3479 n469 VDD GND INV_X1
xU8044 n7438 n870 VDD GND INV_X1
xU8045 n2830 n575 VDD GND INV_X1
xU8046 n2877 n574 VDD GND INV_X1
xU8047 n3061 n573 VDD GND INV_X1
xU8048 n4544 n479 VDD GND INV_X1
xU8049 n1915 n183 VDD GND INV_X1
xU8050 n2677 n217 VDD GND INV_X1
xU8051 n2783 n234 VDD GND INV_X1
xU8052 n2225 n213 VDD GND INV_X1
xU8053 n3891 n293 VDD GND INV_X1
xU8054 n1187 n147 VDD GND INV_X1
xU8055 n4047 n258 VDD GND INV_X1
xU8056 n3116 n198 VDD GND INV_X1
xU8057 n5098 n325 VDD GND INV_X1
xU8058 n3868 n280 VDD GND INV_X1
xU8059 n2249 n224 VDD GND INV_X1
xU8060 n2760 n235 VDD GND INV_X1
xU8061 n1752 n155 VDD GND INV_X1
xU8062 n3000 n205 VDD GND INV_X1
xU8063 n4737 n324 VDD GND INV_X1
xU8064 n4067 n278 VDD GND INV_X1
xU8065 n5319 n315 VDD GND INV_X1
xU8066 n3789 n276 VDD GND INV_X1
xU8067 n3497 n272 VDD GND INV_X1
xU8068 n3990 n283 VDD GND INV_X1
xU8069 n1311 n146 VDD GND INV_X1
xU8070 n4834 n319 VDD GND INV_X1
xU8071 n5464 n347 VDD GND INV_X1
xU8072 n3764 n291 VDD GND INV_X1
xU8073 n2630 n226 VDD GND INV_X1
xU8074 n3694 n271 VDD GND INV_X1
xU8075 n5196 n344 VDD GND INV_X1
xU8076 n5002 n345 VDD GND INV_X1
xU8077 n2810 n210 VDD GND INV_X1
xU8078 n4906 n633 VDD GND INV_X1
xU8079 n3471 n448 VDD GND INV_X1
xU8080 n3671 n295 VDD GND INV_X1
xU8081 n3598 n294 VDD GND INV_X1
xU8082 n2831 n208 VDD GND INV_X1
xU8083 n5297 n316 VDD GND INV_X1
xU8084 n1090 n178 VDD GND INV_X1
xU8085 n2353 n207 VDD GND INV_X1
xU8086 n2852 n223 VDD GND INV_X1
xU8087 n1605 n162 VDD GND INV_X1
xU8088 n1115 n150 VDD GND INV_X1
xU8089 n1504 n142 VDD GND INV_X1
xU8090 n2380 n236 VDD GND INV_X1
xU8091 n5531 n337 VDD GND INV_X1
xU8092 n2979 n204 VDD GND INV_X1
xU8093 n5444 n338 VDD GND INV_X1
xU8094 n1212 n174 VDD GND INV_X1
xU8095 n2438 n212 VDD GND INV_X1
xU8096 n3472 n286 VDD GND INV_X1
xU8097 n4907 n327 VDD GND INV_X1
xU8098 n4091 n292 VDD GND INV_X1
xU8099 n5463 n373 VDD GND INV_X1
xU8100 n4305 n274 VDD GND INV_X1
xU8101 n2326 n202 VDD GND INV_X1
xU8102 n2531 n214 VDD GND INV_X1
xU8103 n4807 n348 VDD GND INV_X1
xU8104 n1310 n527 VDD GND INV_X1
xU8105 n4833 n332 VDD GND INV_X1
xU8106 n2734 n225 VDD GND INV_X1
xU8107 n6808 n850 VDD GND INV_X1
xU8108 n8309 n8290 VDD GND INV_X1
xU8109 n8307 n8287 VDD GND INV_X1
xU8110 n8307 n8286 VDD GND INV_X1
xU8111 n8308 n8289 VDD GND INV_X1
xU8112 n8308 n8288 VDD GND INV_X1
xU8113 n2425 n552 VDD GND INV_X1
xU8114 n5776 n355 VDD GND INV_X1
xU8115 n6823 n848 VDD GND INV_X1
xU8116 n6800 n851 VDD GND INV_X1
xU8117 n2591 n240 VDD GND INV_X1
xU8118 n7014 n836 VDD GND INV_X1
xU8119 n4558 n4570 n4565 VDD GND NAND2_X1
xU8120 n2640 n556 VDD GND INV_X1
xU8121 n7465 n871 VDD GND INV_X1
xU8122 n4550 n482 VDD GND INV_X1
xU8123 n5570 n507 VDD GND INV_X1
xU8124 n5547 n645 n4717 VDD GND NAND2_X1
xU8125 n4278 n4205 n3698 VDD GND NAND2_X1
xU8126 n3297 n562 n2862 VDD GND NAND2_X1
xU8127 n5711 n5712 n5695 VDD GND NOR2_X1
xU8128 n300 n4477 n4461 VDD GND NOR2_X1
xU8129 n4478 n300 VDD GND INV_X1
xU8130 n4276 n619 n3875 VDD GND NAND2_X1
xU8131 n5595 n382 VDD GND INV_X1
xU8132 n2029 n2021 n1858 VDD GND NAND2_X1
xU8133 n3391 n241 n3104 VDD GND NAND2_X1
xU8134 n3153 n431 n3076 VDD GND NAND2_X1
xU8135 n3154 n431 VDD GND INV_X1
xU8136 n7259 n7260 n7217 VDD GND NAND2_X1
xU8137 n3305 n3306 n3087 VDD GND NAND2_X1
xU8138 n3153 n3157 n3150 VDD GND NAND2_X1
xU8139 n3391 n3394 n3389 VDD GND NAND2_X1
xU8140 n2029 n667 n1827 VDD GND NAND2_X1
xU8141 n2025 n667 VDD GND INV_X1
xU8142 n2014 n2020 n1826 VDD GND NAND2_X1
xU8143 n6801 n6802 n6764 VDD GND NAND2_X1
xU8144 n6784 n6764 n6724 VDD GND NAND2_X1
xU8145 n7259 n821 n7243 VDD GND NAND2_X1
xU8146 n7468 n7469 n7410 VDD GND NAND2_X1
xU8147 n3318 n3323 n3086 VDD GND NAND2_X1
xU8148 n4478 n4470 n4458 VDD GND NAND2_X1
xU8149 n7028 n7030 n6996 VDD GND NAND2_X1
xU8150 n5702 n5691 n5503 VDD GND NAND2_X1
xU8151 n5273 n496 VDD GND INV_X1
xU8152 n7474 n7476 n7469 VDD GND NAND2_X1
xU8153 n6811 n6810 n6808 VDD GND NAND2_X1
xU8154 n3648 n451 VDD GND INV_X1
xU8155 n1842 n405 VDD GND INV_X1
xU8156 n1510 n406 VDD GND INV_X1
xU8157 n4720 n640 VDD GND INV_X1
xU8158 n4895 n371 VDD GND INV_X1
xU8159 n2426 n199 VDD GND INV_X1
xU8160 n1515 n399 VDD GND INV_X1
xU8161 n5620 n5621 n5612 VDD GND NAND2_X1
xU8162 n5872 n5867 n5855 VDD GND NAND2_X1
xU8163 n4560 n4564 n4546 VDD GND NAND2_X1
xU8164 n5075 n629 VDD GND INV_X1
xU8165 n3637 n470 VDD GND INV_X1
xU8166 n7483 n7484 n7473 VDD GND NAND2_X1
xU8167 n4384 n4385 n4380 VDD GND NAND2_X1
xU8168 n4886 n342 VDD GND INV_X1
xU8169 n1070 n533 VDD GND INV_X1
xU8170 n3237 n3232 n3227 VDD GND NAND2_X1
xU8171 n2157 n2152 n2140 VDD GND NAND2_X1
xU8172 n4395 n4389 n4377 VDD GND NAND2_X1
xU8173 n2076 n2080 n1917 VDD GND NAND2_X1
xU8174 n1954 n1949 n1937 VDD GND NAND2_X1
xU8175 n1362 n521 VDD GND INV_X1
xU8176 n4468 n4458 n4292 VDD GND NAND2_X1
xU8177 n1129 n148 VDD GND INV_X1
xU8178 n3819 n277 VDD GND INV_X1
xU8179 n1166 n659 VDD GND INV_X1
xU8180 n1852 n182 VDD GND INV_X1
xU8181 n1220 n181 VDD GND INV_X1
xU8182 n3847 n257 VDD GND INV_X1
xU8183 n3856 n474 VDD GND INV_X1
xU8184 n5611 n5612 n5475 VDD GND NAND2_X1
xU8185 n5865 n5855 n5511 VDD GND NAND2_X1
xU8186 n4542 n4546 n4252 VDD GND NAND2_X1
xU8187 n7418 n7373 n7341 VDD GND NAND2_X1
xU8188 n3138 n3227 n3008 VDD GND NAND2_X1
xU8189 n4387 n4377 n4265 VDD GND NAND2_X1
xU8190 n2150 n2140 n1783 VDD GND NAND2_X1
xU8191 n1912 n1917 n1762 VDD GND NAND2_X1
xU8192 n1947 n1937 n1795 VDD GND NAND2_X1
xU8193 n2616 n578 VDD GND INV_X1
xU8194 n4622 n4372 n4284 VDD GND NAND2_X1
xU8195 n1870 n171 VDD GND INV_X1
xU8196 n7217 n7235 n7185 VDD GND NAND2_X1
xU8197 n3308 n3072 n3047 VDD GND NAND2_X1
xU8198 n1604 n173 VDD GND INV_X1
xU8199 n4046 n601 VDD GND INV_X1
xU8200 n1560 n396 VDD GND INV_X1
xU8201 n2653 n227 VDD GND INV_X1
xU8202 n4394 n611 VDD GND INV_X1
xU8203 n1921 n185 VDD GND INV_X1
xU8204 n3243 n581 VDD GND INV_X1
xU8205 n2942 n579 VDD GND INV_X1
xU8206 n5574 n5575 n5415 VDD GND NAND2_X1
xU8207 n3501 n453 VDD GND INV_X1
xU8208 n1102 n530 VDD GND INV_X1
xU8209 n2746 n584 VDD GND INV_X1
xU8210 n1405 n403 VDD GND INV_X1
xU8211 n1021 n663 VDD GND INV_X1
xU8212 n2866 n429 VDD GND INV_X1
xU8213 n1769 n665 VDD GND INV_X1
xU8214 n2261 n585 VDD GND INV_X1
xU8215 n2856 n586 VDD GND INV_X1
xU8216 n1201 n531 VDD GND INV_X1
xU8217 n1114 n657 VDD GND INV_X1
xU8218 n5228 n356 VDD GND INV_X1
xU8219 n990 n658 VDD GND INV_X1
xU8220 n4930 n638 VDD GND INV_X1
xU8221 n2510 n420 VDD GND INV_X1
xU8222 n2608 n419 VDD GND INV_X1
xU8223 n2665 n559 VDD GND INV_X1
xU8224 n1893 n1858 n1774 VDD GND NAND2_X1
xU8225 n3388 n3104 n3030 VDD GND NAND2_X1
xU8226 n3151 n3076 n3039 VDD GND NAND2_X1
xU8227 n6996 n7017 n6962 VDD GND NAND2_X1
xU8228 n3895 n610 VDD GND INV_X1
xU8229 n5218 n502 VDD GND INV_X1
xU8230 n4639 n4632 n4372 VDD GND OR2_X1
xU8231 n4090 n475 VDD GND INV_X1
xU8232 n1785 n158 VDD GND INV_X1
xU8233 n2759 n206 VDD GND INV_X1
xU8234 n5256 n498 VDD GND INV_X1
xU8235 n2248 n555 VDD GND INV_X1
xU8236 n2461 n425 VDD GND INV_X1
xU8237 n5120 n505 VDD GND INV_X1
xU8238 n4015 n604 VDD GND INV_X1
xU8239 n3625 n446 VDD GND INV_X1
xU8240 n2411 n547 VDD GND INV_X1
xU8241 n2999 n576 VDD GND INV_X1
xU8242 n1815 n154 VDD GND INV_X1
xU8243 n2639 n583 VDD GND INV_X1
xU8244 n1336 n157 VDD GND INV_X1
xU8245 n5371 n346 VDD GND INV_X1
xU8246 n4887 n326 VDD GND INV_X1
xU8247 n3820 n263 VDD GND INV_X1
xU8248 n1363 n169 VDD GND INV_X1
xU8249 n2581 n220 VDD GND INV_X1
xU8250 n1816 n139 VDD GND INV_X1
xU8251 n5274 n340 VDD GND INV_X1
xU8252 n3062 n233 VDD GND INV_X1
xU8253 n1561 n144 VDD GND INV_X1
xU8254 n2784 n221 VDD GND INV_X1
xU8255 n5121 n349 VDD GND INV_X1
xU8256 n1167 n170 VDD GND INV_X1
xU8257 n4241 n476 VDD GND INV_X1
xU8258 n4350 n256 VDD GND INV_X1
xU8259 n5076 n341 VDD GND INV_X1
xU8260 n2462 n219 VDD GND INV_X1
xU8261 n4931 n350 VDD GND INV_X1
xU8262 n1382 n152 VDD GND INV_X1
xU8263 n1017 n175 VDD GND INV_X1
xU8264 n3544 n273 VDD GND INV_X1
xU8265 n2412 n200 VDD GND INV_X1
xU8266 n1659 n140 VDD GND INV_X1
xU8267 n2906 n229 VDD GND INV_X1
xU8268 n1871 n138 VDD GND INV_X1
xU8269 n3649 n264 VDD GND INV_X1
xU8270 n2506 n238 VDD GND INV_X1
xU8271 n1258 n165 VDD GND INV_X1
xU8272 n1730 n163 VDD GND INV_X1
xU8273 n2555 n211 VDD GND INV_X1
xU8274 n2678 n230 VDD GND INV_X1
xU8275 n2703 n228 VDD GND INV_X1
xU8276 n3989 n606 VDD GND INV_X1
xU8277 n1284 n177 VDD GND INV_X1
xU8278 n3964 n260 VDD GND INV_X1
xU8279 n5586 n313 VDD GND INV_X1
xU8280 n1532 n149 VDD GND INV_X1
xU8281 n3571 n267 VDD GND INV_X1
xU8282 n1629 n167 VDD GND INV_X1
xU8283 n4782 n329 VDD GND INV_X1
xU8284 n1450 n145 VDD GND INV_X1
xU8285 n2298 n232 VDD GND INV_X1
xU8286 n1503 n401 VDD GND INV_X1
xU8287 n3597 n444 VDD GND INV_X1
xU8288 n1481 n164 VDD GND INV_X1
xU8289 n3934 n288 VDD GND INV_X1
xU8290 n5026 n331 VDD GND INV_X1
xU8291 n3867 n605 VDD GND INV_X1
xU8292 n2437 n423 VDD GND INV_X1
xU8293 n2297 n554 VDD GND INV_X1
xU8294 n4560 n4561 n4552 VDD GND AND2_X1
xU8295 n5872 n5873 n5859 VDD GND AND2_X1
xU8296 n1186 n526 VDD GND INV_X1
xU8297 n1582 n143 VDD GND INV_X1
xU8298 n2352 n553 VDD GND INV_X1
xU8299 n5318 n376 VDD GND INV_X1
xU8300 n4395 n4396 n4381 VDD GND AND2_X1
xU8301 n4465 n4466 n4462 VDD GND AND2_X1
xU8302 n5620 n5624 n5615 VDD GND AND2_X1
xU8303 n2157 n534 n2143 VDD GND AND2_X1
xU8304 n4706 n328 VDD GND INV_X1
xU8305 n5243 n317 VDD GND INV_X1
xU8306 n3848 n279 VDD GND INV_X1
xU8307 n1406 n180 VDD GND INV_X1
xU8308 n3626 n266 VDD GND INV_X1
xU8309 n5049 n318 VDD GND INV_X1
xU8310 n992 n151 VDD GND INV_X1
xU8311 n3788 n284 VDD GND INV_X1
xU8312 n1062 n168 VDD GND INV_X1
xU8313 n5165 n333 VDD GND INV_X1
xU8314 n4016 n275 VDD GND INV_X1
xU8315 n2609 n222 VDD GND INV_X1
xU8316 n4220 n259 VDD GND INV_X1
xU8317 n2554 n422 VDD GND INV_X1
xU8318 n2654 n218 VDD GND INV_X1
xU8319 n1142 n156 VDD GND INV_X1
xU8320 n2799 n239 VDD GND INV_X1
xU8321 n1751 n141 VDD GND INV_X1
xU8322 n5862 n5863 n5858 VDD GND AND2_X1
xU8323 n1351 n532 VDD GND INV_X1
xU8324 n3066 n588 VDD GND INV_X1
xU8325 n5790 n357 VDD GND INV_X1
xU8326 n7027 n834 VDD GND INV_X1
xU8327 n7025 n835 VDD GND INV_X1
xU8328 n2964 n560 VDD GND INV_X1
xU8329 n8340 n8329 VDD GND INV_X1
xU8330 n8340 n8330 VDD GND INV_X1
xU8331 n8340 n8331 VDD GND INV_X1
xU8332 n8281 n8279 VDD GND INV_X1
xU8333 n8281 n8280 VDD GND INV_X1
xU8334 n8281 n8272 VDD GND INV_X1
xU8335 n8281 n8273 VDD GND INV_X1
xU8336 n8281 n8274 VDD GND INV_X1
xU8337 n8281 n8275 VDD GND INV_X1
xU8338 n8281 n8276 VDD GND INV_X1
xU8339 n8281 n8277 VDD GND INV_X1
xU8340 n8281 n8278 VDD GND INV_X1
xU8341 n4942 n506 VDD GND INV_X1
xU8342 n3397 n3398 n3395 VDD GND NAND2_X1
xU8343 n4481 n299 VDD GND INV_X1
xU8344 n1959 n407 VDD GND INV_X1
xU8345 n7054 n837 VDD GND INV_X1
xU8346 n6972 n8247 n8246 VDD GND XOR2_X1
xU8347 n6988 n6989 n8247 VDD GND NAND2_X1
xU8348 n7420 n8249 n8248 VDD GND XOR2_X1
xU8349 n7437 n7438 n8249 VDD GND OR2_X1
xU8350 n7433 n869 VDD GND INV_X1
xU8351 n6749 n849 VDD GND INV_X1
xU8352 n5638 n5628 n5634 VDD GND NAND2_X1
xU8353 n6752 n6753 n6751 VDD GND NAND2_X1
xU8354 n1790 n404 VDD GND INV_X1
xU8355 n5417 n354 VDD GND INV_X1
xU8356 n5414 n5415 n5413 VDD GND NAND2_X1
xU8357 n3510 n285 VDD GND INV_X1
xU8358 n7183 n7238 n7234 VDD GND NAND2_X1
xU8359 n5627 n5628 n5625 VDD GND NAND2_X1
xU8360 n7299 n821 VDD GND INV_X1
xU8361 n7284 n7254 n7271 VDD GND NAND2_X1
xU8362 n6822 n852 VDD GND INV_X1
xU8363 n4631 n457 VDD GND INV_X1
xU8364 n3191 n432 n3161 VDD GND NOR2_X1
xU8365 n3172 n432 VDD GND INV_X1
xU8366 n5817 n5783 n5799 VDD GND NAND2_X1
xU8367 n7304 n822 VDD GND INV_X1
xU8368 n7212 n8250 n7204 VDD GND XOR2_X1
xU8369 n7210 n7211 n8250 VDD GND NAND2_X1
xU8370 n5429 n5486 n4750 VDD GND NAND2_X1
xU8371 n4366 n487 n3511 VDD GND NAND2_X1
xU8372 n4161 n487 VDD GND INV_X1
xU8373 n8326 n5977 n5975 VDD GND NOR2_X1
xU8374 n4324 n4177 n3481 VDD GND NAND2_X1
xU8375 n4620 n4628 n4079 VDD GND NAND2_X1
xU8376 n1840 n1841 n1195 VDD GND NAND2_X1
xU8377 n1786 n2138 n1216 VDD GND NAND2_X1
xU8378 n5991 n8327 n5989 VDD GND NOR2_X1
xU8379 n6131 n8326 n6129 VDD GND NOR2_X1
xU8380 n5984 n8327 n5982 VDD GND NOR2_X1
xU8381 n6033 n8327 n6031 VDD GND NOR2_X1
xU8382 n6145 n8326 n6143 VDD GND NOR2_X1
xU8383 n6075 n8327 n6073 VDD GND NOR2_X1
xU8384 n2147 n2148 n2144 VDD GND NOR2_X1
xU8385 n3123 n3224 n2639 VDD GND NAND2_X1
xU8386 n5492 n5404 n5133 VDD GND NAND2_X1
xU8387 n4318 n4319 n3678 VDD GND NAND2_X1
xU8388 n2194 n2148 n2165 VDD GND NOR2_X1
xU8389 n5591 n5616 n5131 VDD GND NAND2_X1
xU8390 n3083 n3084 n2259 VDD GND NAND2_X1
xU8391 n4355 n4553 n3902 VDD GND NAND2_X1
xU8392 n1931 n1672 n1221 VDD GND NAND2_X1
xU8393 n4333 n4334 n3509 VDD GND NAND2_X1
xU8394 n1876 n1924 n1414 VDD GND NAND2_X1
xU8395 n3175 n3176 n3160 VDD GND NOR2_X1
xU8396 n2936 n435 VDD GND INV_X1
xU8397 n4639 n4640 n4369 VDD GND NOR2_X1
xU8398 n5617 n5618 n5282 VDD GND NAND2_X1
xU8399 n2166 n535 n2154 VDD GND NOR2_X1
xU8400 n2159 n535 VDD GND INV_X1
xU8401 n3088 n3299 n2447 VDD GND NAND2_X1
xU8402 n3017 n246 n2658 VDD GND NAND2_X1
xU8403 n2954 n246 VDD GND INV_X1
xU8404 n3017 n3018 n2619 VDD GND NAND2_X1
xU8405 n4278 n4279 n3659 VDD GND NAND2_X1
xU8406 n3604 n455 VDD GND INV_X1
xU8407 n3098 n3099 n2799 VDD GND NAND2_X1
xU8408 n5771 n5772 n5417 VDD GND NAND2_X1
xU8409 n3023 n2936 n2866 VDD GND NAND2_X1
xU8410 n7252 n7253 n7235 VDD GND NAND2_X1
xU8411 n1837 n1838 n1351 VDD GND NAND2_X1
xU8412 n3318 n3312 n3072 VDD GND NAND2_X1
xU8413 n1904 n1905 n1893 VDD GND NAND2_X1
xU8414 n3400 n3396 n3388 VDD GND NAND2_X1
xU8415 n5562 n363 VDD GND INV_X1
xU8416 n4821 n352 VDD GND INV_X1
xU8417 n1835 n2141 n1648 VDD GND NAND2_X1
xU8418 n4624 n4625 n4193 VDD GND NAND2_X1
xU8419 n4331 n4459 n4131 VDD GND NAND2_X1
xU8420 n3335 n3324 n3308 VDD GND NAND2_X1
xU8421 n5778 n5779 n5575 VDD GND NAND2_X1
xU8422 n7036 n7037 n7025 VDD GND NAND2_X1
xU8423 n6758 n6794 n6654 VDD GND NAND2_X1
xU8424 n5492 n5493 n4720 VDD GND NAND2_X1
xU8425 n7038 n7039 n7014 VDD GND NAND2_X1
xU8426 n3133 n2919 n2856 VDD GND NAND2_X1
xU8427 n7031 n7038 n7017 VDD GND NAND2_X1
xU8428 n2311 n231 VDD GND INV_X1
xU8429 n5805 n358 n5776 VDD GND NAND2_X1
xU8430 n3164 n3172 n3144 VDD GND NAND2_X1
xU8431 n5779 n5783 n5558 VDD GND NAND2_X1
xU8432 n3402 n3403 n3383 VDD GND NAND2_X1
xU8433 n6736 n858 n6637 VDD GND NAND2_X1
xU8434 n6688 n858 VDD GND INV_X1
xU8435 n1072 n402 VDD GND INV_X1
xU8436 n7261 n823 n7239 VDD GND NAND2_X1
xU8437 n1890 n1901 n1769 VDD GND NAND2_X1
xU8438 n3557 n607 VDD GND INV_X1
xU8439 n7252 n7254 n7240 VDD GND NAND2_X1
xU8440 n3335 n3328 n3304 VDD GND NAND2_X1
xU8441 n3021 n564 n3042 VDD GND NAND2_X1
xU8442 n1828 n671 n1225 VDD GND AND2_X1
xU8443 n1687 n671 VDD GND INV_X1
xU8444 n4795 n377 VDD GND INV_X1
xU8445 n1073 n166 VDD GND INV_X1
xU8446 n3400 n3401 n3387 VDD GND NAND2_X1
xU8447 n1904 n666 n1900 VDD GND NAND2_X1
xU8448 n1061 n662 VDD GND INV_X1
xU8449 n5792 n5784 n5574 VDD GND NAND2_X1
xU8450 n4147 n472 VDD GND INV_X1
xU8451 n7189 n7151 n7212 VDD GND NAND2_X1
xU8452 n4771 n335 VDD GND INV_X1
xU8453 n3530 n449 VDD GND INV_X1
xU8454 n5486 n5487 n5086 VDD GND AND2_X1
xU8455 n2965 n3088 n2665 VDD GND NAND2_X1
xU8456 n5164 n504 VDD GND INV_X1
xU8457 n2313 n577 VDD GND INV_X1
xU8458 n6824 n6805 n6784 VDD GND NAND2_X1
xU8459 n4366 n4367 n4056 VDD GND AND2_X1
xU8460 n3739 n290 VDD GND INV_X1
xU8461 n4457 n4458 n4204 VDD GND NAND2_X1
xU8462 n428 n3158 n3151 VDD GND NAND2_X1
xU8463 n3168 n428 VDD GND INV_X1
xU8464 n5617 n5384 n5595 VDD GND NAND2_X1
xU8465 n7475 n7469 n7374 VDD GND NAND2_X1
xU8466 n5619 n5612 n5383 VDD GND NAND2_X1
xU8467 n5854 n5855 n5403 VDD GND NAND2_X1
xU8468 n4543 n4546 n4160 VDD GND NAND2_X1
xU8469 n4376 n4377 n4186 VDD GND NAND2_X1
xU8470 n1913 n1917 n1671 VDD GND NAND2_X1
xU8471 n5774 n5575 n5517 VDD GND NAND2_X1
xU8472 n7017 n6997 n6964 VDD GND NAND2_X1
xU8473 n3151 n3077 n3036 VDD GND NAND2_X1
xU8474 n3388 n3105 n3032 VDD GND NAND2_X1
xU8475 n1893 n1859 n1775 VDD GND NAND2_X1
xU8476 n1918 n1919 n1912 VDD GND NAND2_X1
xU8477 n4397 n4401 n4387 VDD GND NAND2_X1
xU8478 n3240 n3241 n3138 VDD GND NAND2_X1
xU8479 n4547 n4548 n4542 VDD GND NAND2_X1
xU8480 n4507 n304 VDD GND INV_X1
xU8481 n4976 n636 VDD GND INV_X1
xU8482 n1257 n528 VDD GND INV_X1
xU8483 n5205 n375 VDD GND INV_X1
xU8484 n5690 n5691 n5428 VDD GND NAND2_X1
xU8485 n4371 n4372 n4176 VDD GND NAND2_X1
xU8486 n5611 n5619 n5477 VDD GND NAND2_X1
xU8487 n1947 n1936 n1792 VDD GND NAND2_X1
xU8488 n1912 n1913 n1764 VDD GND NAND2_X1
xU8489 n5865 n5854 n5508 VDD GND NAND2_X1
xU8490 n4387 n4376 n4267 VDD GND NAND2_X1
xU8491 n3138 n3139 n3010 VDD GND NAND2_X1
xU8492 n4622 n4371 n4286 VDD GND NAND2_X1
xU8493 n4542 n4543 n4254 VDD GND NAND2_X1
xU8494 n4468 n4457 n4293 VDD GND NAND2_X1
xU8495 n7468 n7475 n7412 VDD GND NAND2_X1
xU8496 n1799 n1697 n1842 VDD GND NAND2_X1
xU8497 n1799 n1800 n1510 VDD GND NAND2_X1
xU8498 n4020 n612 VDD GND INV_X1
xU8499 n2138 n540 VDD GND INV_X1
xU8500 n2150 n2139 n1780 VDD GND NAND2_X1
xU8501 n5605 n5775 n5419 VDD GND NAND2_X1
xU8502 n1896 n1897 n1703 VDD GND NAND2_X1
xU8503 n4562 n4563 n4554 VDD GND NAND2_X1
xU8504 n3229 n3231 n3226 VDD GND NAND2_X1
xU8505 n2078 n2079 n1925 VDD GND NAND2_X1
xU8506 n3795 n297 VDD GND INV_X1
xU8507 n5709 n5717 n5702 VDD GND NAND2_X1
xU8508 n7189 n7190 n7108 VDD GND NAND2_X1
xU8509 n5632 n5626 n5611 VDD GND NAND2_X1
xU8510 n1956 n1960 n1947 VDD GND NAND2_X1
xU8511 n4475 n4482 n4468 VDD GND NAND2_X1
xU8512 n5874 n5880 n5865 VDD GND NAND2_X1
xU8513 n2158 n2163 n2150 VDD GND NAND2_X1
xU8514 n4637 n458 n4622 VDD GND NAND2_X1
xU8515 n4644 n458 VDD GND INV_X1
xU8516 n7481 n7477 n7468 VDD GND NAND2_X1
xU8517 n4591 n4555 n4570 VDD GND NAND2_X1
xU8518 n4576 n484 VDD GND INV_X1
xU8519 n5882 n5875 n5869 VDD GND NAND2_X1
xU8520 n5886 n644 VDD GND INV_X1
xU8521 n6792 n859 n6720 VDD GND NAND2_X1
xU8522 n5692 n514 n5498 VDD GND NAND2_X1
xU8523 n4315 n623 n4033 VDD GND NAND2_X1
xU8524 n4272 n461 n4280 VDD GND NAND2_X1
xU8525 n4374 n620 n4261 VDD GND NAND2_X1
xU8526 n4455 n305 n4288 VDD GND NAND2_X1
xU8527 n4357 n488 n4248 VDD GND NAND2_X1
xU8528 n7461 n877 n7406 VDD GND NAND2_X1
xU8529 n3379 n247 n3026 VDD GND NAND2_X1
xU8530 n7439 n881 n7420 VDD GND NAND2_X1
xU8531 n6970 n6931 n6897 VDD GND NAND2_X1
xU8532 n3079 n438 n2594 VDD GND NAND2_X1
xU8533 n3308 n3073 n3044 VDD GND NAND2_X1
xU8534 n7214 n7242 n7221 VDD GND NAND2_X1
xU8535 n1894 n675 n1614 VDD GND NAND2_X1
xU8536 n4397 n614 n4383 VDD GND NAND2_X1
xU8537 n4547 n4555 n4551 VDD GND NAND2_X1
xU8538 n1918 n1926 n1922 VDD GND NAND2_X1
xU8539 n3240 n3248 n3225 VDD GND NAND2_X1
xU8540 n7474 n873 n7466 VDD GND NAND2_X1
xU8541 n1936 n1937 n1696 VDD GND NAND2_X1
xU8542 n2139 n2140 n1715 VDD GND NAND2_X1
xU8543 n5702 n5690 n5500 VDD GND NAND2_X1
xU8544 n3081 n3155 n2894 VDD GND NAND2_X1
xU8545 n3096 n3392 n2890 VDD GND NAND2_X1
xU8546 n5519 n5520 n5412 VDD GND NAND2_X1
xU8547 n2031 n670 VDD GND INV_X1
xU8548 n482 n4362 n4124 VDD GND NAND2_X1
xU8549 n6993 n7012 n7000 VDD GND NAND2_X1
xU8550 n185 n1881 n1636 VDD GND NAND2_X1
xU8551 n581 n3129 n2884 VDD GND NAND2_X1
xU8552 n5791 n5792 n5559 VDD GND AND2_X1
xU8553 n6801 n6803 n6796 VDD GND AND2_X1
xU8554 n7028 n7029 n7013 VDD GND AND2_X1
xU8555 n4187 n619 VDD GND INV_X1
xU8556 n3374 n562 VDD GND INV_X1
xU8557 n5571 n5572 n4939 VDD GND AND2_X1
xU8558 n4032 n608 VDD GND INV_X1
xU8559 n3171 n3309 n2967 VDD GND NAND2_X1
xU8560 n508 n5704 n5691 VDD GND NAND2_X1
xU8561 n5711 n508 VDD GND INV_X1
xU8562 n6996 n6997 n6930 VDD GND NAND2_X1
xU8563 n1858 n1859 n1686 VDD GND NAND2_X1
xU8564 n3104 n3105 n2953 VDD GND NAND2_X1
xU8565 n7218 n7235 n7183 VDD GND NAND2_X1
xU8566 n871 n7463 n7353 VDD GND NAND2_X1
xU8567 n6824 n6815 n6785 VDD GND AND2_X1
xU8568 n5852 n649 n5506 VDD GND NAND2_X1
xU8569 n3072 n3073 n2964 VDD GND NAND2_X1
xU8570 n3076 n3077 n2935 VDD GND NAND2_X1
xU8571 n6763 n6764 n6687 VDD GND NAND2_X1
xU8572 n611 n4378 n4136 VDD GND NAND2_X1
xU8573 n4749 n635 VDD GND INV_X1
xU8574 n1792 n1946 n1700 VDD GND NAND2_X1
xU8575 n4004 n445 VDD GND INV_X1
xU8576 n4293 n4467 n4208 VDD GND NAND2_X1
xU8577 n3032 n3384 n2957 VDD GND NAND2_X1
xU8578 n5508 n5864 n5407 VDD GND NAND2_X1
xU8579 n5477 n5599 n5387 VDD GND NAND2_X1
xU8580 n3428 n3403 n3397 VDD GND NAND2_X1
xU8581 n2060 n2020 n1909 VDD GND NAND2_X1
xU8582 n3586 n456 VDD GND INV_X1
xU8583 n5639 n383 n5628 VDD GND NAND2_X1
xU8584 n6784 n6763 n6726 VDD GND NAND2_X1
xU8585 n5927 n645 VDD GND INV_X1
xU8586 n2045 n666 n2023 VDD GND NAND2_X1
xU8587 n3139 n3227 n3066 VDD GND NAND2_X1
xU8588 n4571 n4563 n4558 VDD GND NAND2_X1
xU8589 n4253 n486 VDD GND INV_X1
xU8590 n4128 n452 VDD GND INV_X1
xU8591 n874 n7484 n7480 VDD GND NAND2_X1
xU8592 n7526 n874 VDD GND INV_X1
xU8593 n3168 n3176 n3152 VDD GND OR2_X1
xU8594 n4101 n609 VDD GND INV_X1
xU8595 n6850 n6811 n6806 VDD GND NAND2_X1
xU8596 n5517 n5777 n5183 VDD GND NAND2_X1
xU8597 n4254 n4359 n4164 VDD GND NAND2_X1
xU8598 n7067 n7037 n7034 VDD GND NAND2_X1
xU8599 n7076 n838 VDD GND INV_X1
xU8600 n3276 n3231 n3246 VDD GND NAND2_X1
xU8601 n3287 n589 VDD GND INV_X1
xU8602 n2083 n2079 n1929 VDD GND NAND2_X1
xU8603 n2090 n187 VDD GND INV_X1
xU8604 n4035 n298 VDD GND INV_X1
xU8605 n4433 n4385 n4403 VDD GND NAND2_X1
xU8606 n4444 n616 VDD GND INV_X1
xU8607 n7217 n7218 n7150 VDD GND NAND2_X1
xU8608 n4675 n4630 n4646 VDD GND NAND2_X1
xU8609 n4517 n4465 n4484 VDD GND NAND2_X1
xU8610 n5664 n5631 n5627 VDD GND NAND2_X1
xU8611 n2416 n558 VDD GND INV_X1
xU8612 n5774 n5574 n5519 VDD GND NAND2_X1
xU8613 n7272 n823 n7258 VDD GND NAND2_X1
xU8614 n5747 n5700 n5719 VDD GND NAND2_X1
xU8615 n1992 n1945 n1962 VDD GND NAND2_X1
xU8616 n5485 n503 VDD GND INV_X1
xU8617 n3903 n480 VDD GND INV_X1
xU8618 n5545 n637 VDD GND INV_X1
xU8619 n3074 n427 VDD GND INV_X1
xU8620 n1829 n529 VDD GND INV_X1
xU8621 n4404 n614 n4391 VDD GND NAND2_X1
xU8622 n5726 n512 VDD GND INV_X1
xU8623 n4736 n351 VDD GND INV_X1
xU8624 n2273 n216 VDD GND INV_X1
xU8625 n5342 n339 VDD GND INV_X1
xU8626 n4117 n268 VDD GND INV_X1
xU8627 n2878 n215 VDD GND INV_X1
xU8628 n4977 n334 VDD GND INV_X1
xU8629 n4707 n353 VDD GND INV_X1
xU8630 n1429 n176 VDD GND INV_X1
xU8631 n5144 n321 VDD GND INV_X1
xU8632 n1041 n160 VDD GND INV_X1
xU8633 n3522 n261 VDD GND INV_X1
xU8634 n3718 n289 VDD GND INV_X1
xU8635 n4761 n336 VDD GND INV_X1
xU8636 n4953 n322 VDD GND INV_X1
xU8637 n4148 n287 VDD GND INV_X1
xU8638 n1236 n159 VDD GND INV_X1
xU8639 n3740 n265 VDD GND INV_X1
xU8640 n3914 n270 VDD GND INV_X1
xU8641 n5630 n5631 n5623 VDD GND AND2_X1
xU8642 n5709 n5710 n5698 VDD GND AND2_X1
xU8643 n7481 n7482 n7467 VDD GND AND2_X1
xU8644 n4637 n4638 n4629 VDD GND AND2_X1
xU8645 n4475 n4476 n4464 VDD GND AND2_X1
xU8646 n3237 n3244 n3230 VDD GND AND2_X1
xU8647 n1954 n1955 n1941 VDD GND AND2_X1
xU8648 n2076 n2077 n1923 VDD GND AND2_X1
xU8649 n5500 n5701 n5433 VDD GND AND2_X1
xU8650 n3044 n3310 n2721 VDD GND AND2_X1
xU8651 n5699 n5700 n5696 VDD GND AND2_X1
xU8652 n1944 n1945 n1940 VDD GND AND2_X1
xU8653 n5874 n5875 n5861 VDD GND AND2_X1
xU8654 n4862 n314 VDD GND INV_X1
xU8655 n2483 n201 VDD GND INV_X1
xU8656 n457 n4630 n4370 VDD GND AND2_X1
xU8657 n4329 n308 n3834 VDD GND AND2_X1
xU8658 n1803 n672 n1770 VDD GND AND2_X1
xU8659 n3417 n241 VDD GND INV_X1
xU8660 n5632 n383 n5614 VDD GND AND2_X1
xU8661 n2158 n2159 n2146 VDD GND AND2_X1
xU8662 n1956 n1957 n1943 VDD GND AND2_X1
xU8663 n3094 n250 n2798 VDD GND AND2_X1
xU8664 n2181 n534 VDD GND INV_X1
xU8665 n3438 n244 VDD GND INV_X1
xU8666 n3978 n477 VDD GND INV_X1
xU8667 n6019 n8335 n6017 VDD GND AND2_X1
xU8668 n6089 n8334 n6087 VDD GND AND2_X1
xU8669 n8339 n5963 n5961 VDD GND AND2_X1
xU8670 n5881 n5869 n5879 VDD GND NAND2_X1
xU8671 n6806 n6807 n6804 VDD GND NAND2_X1
xU8672 n1909 n2023 n2040 VDD GND NAND2_X1
xU8673 n8245 n8340 VDD GND BUF_X1
xU8674 n8401 n8431 VDD GND BUF_X1
xU8675 n8401 n8429 VDD GND BUF_X1
xU8676 n8401 n8432 VDD GND BUF_X1
xU8677 n8401 n8430 VDD GND BUF_X1
xU8678 n8401 n8428 VDD GND BUF_X1
xU8679 n8377 n8396 VDD GND BUF_X1
xU8680 n8377 n8397 VDD GND BUF_X1
xU8681 n8375 n8392 VDD GND BUF_X1
xU8682 n8376 n8394 VDD GND BUF_X1
xU8683 n8374 n8389 VDD GND BUF_X1
xU8684 n8376 n8395 VDD GND BUF_X1
xU8685 n8376 n8393 VDD GND BUF_X1
xU8686 n8375 n8390 VDD GND BUF_X1
xU8687 n8375 n8391 VDD GND BUF_X1
xU8688 n8400 n8423 VDD GND BUF_X1
xU8689 n8374 n8388 VDD GND BUF_X1
xU8690 n1009 n8348 VDD GND BUF_X1
xU8691 n1009 n8347 VDD GND BUF_X1
xU8692 n1009 n8350 VDD GND BUF_X1
xU8693 n1009 n8346 VDD GND BUF_X1
xU8694 n1009 n8349 VDD GND BUF_X1
xU8695 n8399 n8411 VDD GND BUF_X1
xU8696 n8399 n8408 VDD GND BUF_X1
xU8697 n8399 n8410 VDD GND BUF_X1
xU8698 n8399 n8409 VDD GND BUF_X1
xU8699 n8400 n8422 VDD GND BUF_X1
xU8700 n8400 n8419 VDD GND BUF_X1
xU8701 n8400 n8421 VDD GND BUF_X1
xU8702 n8400 n8420 VDD GND BUF_X1
xU8703 n8399 n8412 VDD GND BUF_X1
xU8704 n8374 n8387 VDD GND BUF_X1
xU8705 n8372 n8381 VDD GND BUF_X1
xU8706 n8371 n8379 VDD GND BUF_X1
xU8707 n8371 n8378 VDD GND BUF_X1
xU8708 n8372 n8382 VDD GND BUF_X1
xU8709 n8373 n8386 VDD GND BUF_X1
xU8710 n8373 n8385 VDD GND BUF_X1
xU8711 n8372 n8383 VDD GND BUF_X1
xU8712 n8373 n8384 VDD GND BUF_X1
xU8713 n8371 n8380 VDD GND BUF_X1
xU8714 n8310 n8313 VDD GND BUF_X1
xU8715 n8354 n8364 VDD GND BUF_X1
xU8716 n8355 n8368 VDD GND BUF_X1
xU8717 n8354 n8363 VDD GND BUF_X1
xU8718 n8355 n8366 VDD GND BUF_X1
xU8719 n8353 n8361 VDD GND BUF_X1
xU8720 n8355 n8367 VDD GND BUF_X1
xU8721 n8354 n8365 VDD GND BUF_X1
xU8722 n8353 n8362 VDD GND BUF_X1
xU8723 n8310 n8315 VDD GND BUF_X1
xU8724 n8310 n8317 VDD GND BUF_X1
xU8725 n8310 n8314 VDD GND BUF_X1
xU8726 n8311 n8318 VDD GND BUF_X1
xU8727 n8310 n8316 VDD GND BUF_X1
xU8728 n8311 n8319 VDD GND BUF_X1
xU8729 n8311 n8322 VDD GND BUF_X1
xU8730 n8311 n8320 VDD GND BUF_X1
xU8731 n8311 n8321 VDD GND BUF_X1
xU8732 n8312 n8323 VDD GND BUF_X1
xU8733 n8312 n8324 VDD GND BUF_X1
xU8734 n8356 n8369 VDD GND BUF_X1
xU8735 n8312 n8325 VDD GND BUF_X1
xU8736 n8255 n8258 VDD GND BUF_X1
xU8737 n8256 n8267 VDD GND BUF_X1
xU8738 n8256 n8266 VDD GND BUF_X1
xU8739 n8256 n8265 VDD GND BUF_X1
xU8740 n8256 n8263 VDD GND BUF_X1
xU8741 n8255 n8262 VDD GND BUF_X1
xU8742 n8255 n8261 VDD GND BUF_X1
xU8743 n8255 n8260 VDD GND BUF_X1
xU8744 n8255 n8259 VDD GND BUF_X1
xU8745 n8256 n8264 VDD GND BUF_X1
xU8746 n8257 n8270 VDD GND BUF_X1
xU8747 n8257 n8269 VDD GND BUF_X1
xU8748 n8257 n8268 VDD GND BUF_X1
xU8749 n8353 n8360 VDD GND BUF_X1
xU8750 n8352 n8357 VDD GND BUF_X1
xU8751 n8352 n8358 VDD GND BUF_X1
xU8752 n8352 n8359 VDD GND BUF_X1
xU8753 n8245 n8338 VDD GND BUF_X1
xU8754 n8245 n8335 VDD GND BUF_X1
xU8755 n8245 n8336 VDD GND BUF_X1
xU8756 n8245 n8337 VDD GND BUF_X1
xU8757 n8245 n8339 VDD GND BUF_X1
xU8758 n8338 n8333 VDD GND BUF_X1
xU8759 n8336 n8332 VDD GND BUF_X1
xU8760 n8339 n8334 VDD GND BUF_X1
xU8761 n6610 n8282 VDD GND BUF_X1
xU8762 n6610 n8283 VDD GND BUF_X1
xU8763 n6610 n8284 VDD GND BUF_X1
xU8764 n6610 n8285 VDD GND BUF_X1
xU8765 n5500 n5501 n5499 VDD GND NAND2_X1
xU8766 n4254 n4255 n4250 VDD GND NAND2_X1
xU8767 n1764 n1765 n1760 VDD GND NAND2_X1
xU8768 n3032 n3033 n3028 VDD GND NAND2_X1
xU8769 n3036 n3037 n3035 VDD GND NAND2_X1
xU8770 n5477 n5478 n5473 VDD GND NAND2_X1
xU8771 n4286 n4287 n4282 VDD GND NAND2_X1
xU8772 n3010 n3011 n3006 VDD GND NAND2_X1
xU8773 n1792 n1793 n1791 VDD GND NAND2_X1
xU8774 n5508 n5509 n5507 VDD GND NAND2_X1
xU8775 n1775 n1776 n1772 VDD GND NAND2_X1
xU8776 n7207 n7246 n7241 VDD GND AND2_X1
xU8777 n5821 n360 VDD GND INV_X1
xU8778 n2196 n537 VDD GND INV_X1
xU8779 n6765 n6766 n6760 VDD GND NAND2_X1
xU8780 n4267 n4268 n4263 VDD GND NAND2_X1
xU8781 n4293 n4294 n4290 VDD GND NAND2_X1
xU8782 n5667 n384 VDD GND INV_X1
xU8783 n7211 n7215 n7233 VDD GND NAND2_X1
xU8784 n4500 n302 VDD GND INV_X1
xU8785 n5673 n387 VDD GND INV_X1
xU8786 n6834 n855 VDD GND INV_X1
xU8787 n6756 n862 n6754 VDD GND NAND2_X1
xU8788 n7182 n820 n7181 VDD GND NOR2_X1
xU8789 n7183 n820 VDD GND INV_X1
xU8790 n7412 n7413 n7408 VDD GND NAND2_X1
xU8791 n6752 n6759 n6782 VDD GND NAND2_X1
xU8792 n6726 n6727 n6722 VDD GND NAND2_X1
xU8793 n6964 n6965 n6960 VDD GND NAND2_X1
xU8794 n870 n7441 n7470 VDD GND NAND2_X1
xU8795 n6989 n6994 n7022 VDD GND NAND2_X1
xU8796 n6929 n6930 n6926 VDD GND NAND2_X1
xU8797 n5901 n641 VDD GND INV_X1
xU8798 n1984 n408 VDD GND INV_X1
xU8799 n7277 n823 VDD GND INV_X1
xU8800 n5703 n510 VDD GND INV_X1
xU8801 n1780 n1781 n1779 VDD GND NAND2_X1
xU8802 n3044 n569 n3043 VDD GND NAND2_X1
xU8803 n3045 n569 VDD GND INV_X1
xU8804 n5517 n5518 n5516 VDD GND NAND2_X1
xU8805 n5640 n383 VDD GND INV_X1
xU8806 n7149 n7150 n7146 VDD GND NAND2_X1
xU8807 n3327 n3328 n3314 VDD GND AND2_X1
xU8808 n3415 n242 VDD GND INV_X1
xU8809 n6817 n853 VDD GND INV_X1
xU8810 n3083 n3082 n2308 VDD GND NAND2_X1
xU8811 n3297 n3298 n2416 VDD GND NAND2_X1
xU8812 n6138 n8326 n6136 VDD GND NOR2_X1
xU8813 n8328 n6327 n6325 VDD GND NOR2_X1
xU8814 n8327 n6271 n6269 VDD GND NOR2_X1
xU8815 n8327 n6159 n6157 VDD GND NOR2_X1
xU8816 n8328 n6383 n6381 VDD GND NOR2_X1
xU8817 n8328 n6320 n6318 VDD GND NOR2_X1
xU8818 n8327 n6264 n6262 VDD GND NOR2_X1
xU8819 n8327 n6152 n6150 VDD GND NOR2_X1
xU8820 n8328 n6376 n6374 VDD GND NOR2_X1
xU8821 n8327 n6187 n6185 VDD GND NOR2_X1
xU8822 n8327 n6124 n6122 VDD GND NOR2_X1
xU8823 n8328 n6348 n6346 VDD GND NOR2_X1
xU8824 n8327 n6285 n6283 VDD GND NOR2_X1
xU8825 n8327 n6229 n6227 VDD GND NOR2_X1
xU8826 n8327 n6201 n6199 VDD GND NOR2_X1
xU8827 n8327 n6236 n6234 VDD GND NOR2_X1
xU8828 n8327 n6173 n6171 VDD GND NOR2_X1
xU8829 n8328 n6341 n6339 VDD GND NOR2_X1
xU8830 n8328 n6397 n6395 VDD GND NOR2_X1
xU8831 n8328 n6460 n6458 VDD GND NOR2_X1
xU8832 n8328 n6425 n6423 VDD GND NOR2_X1
xU8833 n8328 n6453 n6451 VDD GND NOR2_X1
xU8834 n8327 n6292 n6290 VDD GND NOR2_X1
xU8835 n8328 n6411 n6409 VDD GND NOR2_X1
xU8836 n8327 n6194 n6192 VDD GND NOR2_X1
xU8837 n8328 n6418 n6416 VDD GND NOR2_X1
xU8838 n8326 n6103 n6101 VDD GND NOR2_X1
xU8839 n8326 n6047 n6045 VDD GND NOR2_X1
xU8840 n8326 n6040 n6038 VDD GND NOR2_X1
xU8841 n8326 n6012 n6010 VDD GND NOR2_X1
xU8842 n8326 n6068 n6066 VDD GND NOR2_X1
xU8843 n8326 n5970 n5968 VDD GND NOR2_X1
xU8844 n5561 n5607 n4711 VDD GND NAND2_X1
xU8845 n3023 n3024 n2369 VDD GND NAND2_X1
xU8846 n1931 n2075 n1394 VDD GND NAND2_X1
xU8847 n1671 n1820 n1540 VDD GND NAND2_X1
xU8848 n4276 n4277 n3801 VDD GND NAND2_X1
xU8849 n1786 n1787 n1004 VDD GND NAND2_X1
xU8850 n5488 n5489 n5410 VDD GND NOR2_X1
xU8851 n6026 n8326 n6024 VDD GND NOR2_X1
xU8852 n6082 n8327 n6080 VDD GND NOR2_X1
xU8853 n5940 n8326 n5938 VDD GND NOR2_X1
xU8854 n6054 n8326 n6052 VDD GND NOR2_X1
xU8855 n6110 n8327 n6108 VDD GND NOR2_X1
xU8856 n5733 n5712 n5707 VDD GND NOR2_X1
xU8857 n3133 n3134 n2819 VDD GND NAND2_X1
xU8858 n5771 n5782 n5326 VDD GND NAND2_X1
xU8859 n3145 n3146 n2595 VDD GND NAND2_X1
xU8860 n4176 n4326 n3586 VDD GND NAND2_X1
xU8861 n5777 n5840 n5822 VDD GND NAND2_X1
xU8862 n5490 n5773 n5515 VDD GND NAND2_X1
xU8863 n5513 n652 VDD GND INV_X1
xU8864 n3066 n3067 n2748 VDD GND NAND2_X1
xU8865 n5728 n514 VDD GND INV_X1
xU8866 n6860 n863 VDD GND INV_X1
xU8867 n3333 n564 VDD GND INV_X1
xU8868 n5805 n5797 n5774 VDD GND NAND2_X1
xU8869 n1828 n2012 n1197 VDD GND NAND2_X1
xU8870 n3375 n567 VDD GND INV_X1
xU8871 n5552 n5856 n5355 VDD GND NAND2_X1
xU8872 n7459 n7460 n7379 VDD GND NAND2_X1
xU8873 n5597 n5598 n5348 VDD GND NAND2_X1
xU8874 n1847 n1938 n1643 VDD GND NAND2_X1
xU8875 n5568 n5693 n5360 VDD GND NAND2_X1
xU8876 n7040 n7036 n6997 VDD GND NAND2_X1
xU8877 n1906 n2014 n1859 VDD GND NAND2_X1
xU8878 n3311 n3305 n3073 VDD GND NAND2_X1
xU8879 n3163 n3164 n3077 VDD GND NAND2_X1
xU8880 n3123 n3124 n2915 VDD GND NAND2_X1
xU8881 n1933 n1934 n1790 VDD GND NAND2_X1
xU8882 n3404 n3402 n3105 VDD GND NAND2_X1
xU8883 n4620 n4621 n4171 VDD GND NAND2_X1
xU8884 n4333 n4332 n4199 VDD GND NAND2_X1
xU8885 n5591 n5592 n5378 VDD GND NAND2_X1
xU8886 n5547 n5553 n5398 VDD GND NAND2_X1
xU8887 n1837 n1836 n1710 VDD GND NAND2_X1
xU8888 n1840 n1848 n1691 VDD GND NAND2_X1
xU8889 n1876 n1877 n1666 VDD GND NAND2_X1
xU8890 n4355 n4356 n4155 VDD GND NAND2_X1
xU8891 n3098 n3097 n2948 VDD GND NAND2_X1
xU8892 n7255 n7261 n7218 VDD GND NAND2_X1
xU8893 n6809 n6810 n6763 VDD GND NAND2_X1
xU8894 n7244 n7250 n7191 VDD GND NAND2_X1
xU8895 n4467 n4523 n4504 VDD GND NAND2_X1
xU8896 n3121 n3122 n3004 VDD GND NAND2_X1
xU8897 n2004 n414 VDD GND INV_X1
xU8898 n1696 n1839 n1299 VDD GND AND2_X1
xU8899 n1878 n1879 n1758 VDD GND NAND2_X1
xU8900 n2135 n2136 n1778 VDD GND NAND2_X1
xU8901 n7015 n7035 n6958 VDD GND NAND2_X1
xU8902 n5593 n5594 n5471 VDD GND NAND2_X1
xU8903 n5889 n649 VDD GND INV_X1
xU8904 n6134 n6135 n8002 VDD GND NAND2_X1
xU8905 n6139 n6140 n6134 VDD GND NOR2_X1
xU8906 n6136 n6137 n6135 VDD GND NOR2_X1
xU8907 n8315 n29 n6139 VDD GND NOR2_X1
xU8908 n6323 n6324 n8029 VDD GND NAND2_X1
xU8909 n6328 n6329 n6323 VDD GND NOR2_X1
xU8910 n6325 n6326 n6324 VDD GND NOR2_X1
xU8911 n8318 n56 n6328 VDD GND NOR2_X1
xU8912 n6267 n6268 n8021 VDD GND NAND2_X1
xU8913 n6272 n6273 n6267 VDD GND NOR2_X1
xU8914 n6269 n6270 n6268 VDD GND NOR2_X1
xU8915 n8317 n48 n6272 VDD GND NOR2_X1
xU8916 n6155 n6156 n8005 VDD GND NAND2_X1
xU8917 n6160 n6161 n6155 VDD GND NOR2_X1
xU8918 n6157 n6158 n6156 VDD GND NOR2_X1
xU8919 n8316 n32 n6160 VDD GND NOR2_X1
xU8920 n6379 n6380 n8037 VDD GND NAND2_X1
xU8921 n6384 n6385 n6379 VDD GND NOR2_X1
xU8922 n6381 n6382 n6380 VDD GND NOR2_X1
xU8923 n8319 n64 n6384 VDD GND NOR2_X1
xU8924 n6316 n6317 n8028 VDD GND NAND2_X1
xU8925 n6321 n6322 n6316 VDD GND NOR2_X1
xU8926 n6318 n6319 n6317 VDD GND NOR2_X1
xU8927 n8318 n55 n6321 VDD GND NOR2_X1
xU8928 n6260 n6261 n8020 VDD GND NAND2_X1
xU8929 n6265 n6266 n6260 VDD GND NOR2_X1
xU8930 n6262 n6263 n6261 VDD GND NOR2_X1
xU8931 n8317 n47 n6265 VDD GND NOR2_X1
xU8932 n6148 n6149 n8004 VDD GND NAND2_X1
xU8933 n6153 n6154 n6148 VDD GND NOR2_X1
xU8934 n6150 n6151 n6149 VDD GND NOR2_X1
xU8935 n8316 n31 n6153 VDD GND NOR2_X1
xU8936 n6372 n6373 n8036 VDD GND NAND2_X1
xU8937 n6377 n6378 n6372 VDD GND NOR2_X1
xU8938 n6374 n6375 n6373 VDD GND NOR2_X1
xU8939 n8319 n63 n6377 VDD GND NOR2_X1
xU8940 n6183 n6184 n8009 VDD GND NAND2_X1
xU8941 n6188 n6189 n6183 VDD GND NOR2_X1
xU8942 n6185 n6186 n6184 VDD GND NOR2_X1
xU8943 n8316 n36 n6188 VDD GND NOR2_X1
xU8944 n6120 n6121 n8000 VDD GND NAND2_X1
xU8945 n6125 n6126 n6120 VDD GND NOR2_X1
xU8946 n6122 n6123 n6121 VDD GND NOR2_X1
xU8947 n8315 n27 n6125 VDD GND NOR2_X1
xU8948 n6344 n6345 n8032 VDD GND NAND2_X1
xU8949 n6349 n6350 n6344 VDD GND NOR2_X1
xU8950 n6346 n6347 n6345 VDD GND NOR2_X1
xU8951 n8318 n59 n6349 VDD GND NOR2_X1
xU8952 n6281 n6282 n8023 VDD GND NAND2_X1
xU8953 n6286 n6287 n6281 VDD GND NOR2_X1
xU8954 n6283 n6284 n6282 VDD GND NOR2_X1
xU8955 n8317 n50 n6286 VDD GND NOR2_X1
xU8956 n6225 n6226 n8015 VDD GND NAND2_X1
xU8957 n6230 n6231 n6225 VDD GND NOR2_X1
xU8958 n6227 n6228 n6226 VDD GND NOR2_X1
xU8959 n8317 n42 n6230 VDD GND NOR2_X1
xU8960 n6197 n6198 n8011 VDD GND NAND2_X1
xU8961 n6202 n6203 n6197 VDD GND NOR2_X1
xU8962 n6199 n6200 n6198 VDD GND NOR2_X1
xU8963 n8316 n38 n6202 VDD GND NOR2_X1
xU8964 n6232 n6233 n8016 VDD GND NAND2_X1
xU8965 n6237 n6238 n6232 VDD GND NOR2_X1
xU8966 n6234 n6235 n6233 VDD GND NOR2_X1
xU8967 n8317 n43 n6237 VDD GND NOR2_X1
xU8968 n6169 n6170 n8007 VDD GND NAND2_X1
xU8969 n6174 n6175 n6169 VDD GND NOR2_X1
xU8970 n6171 n6172 n6170 VDD GND NOR2_X1
xU8971 n8316 n34 n6174 VDD GND NOR2_X1
xU8972 n6337 n6338 n8031 VDD GND NAND2_X1
xU8973 n6342 n6343 n6337 VDD GND NOR2_X1
xU8974 n6339 n6340 n6338 VDD GND NOR2_X1
xU8975 n8318 n58 n6342 VDD GND NOR2_X1
xU8976 n6393 n6394 n8039 VDD GND NAND2_X1
xU8977 n6398 n6399 n6393 VDD GND NOR2_X1
xU8978 n6395 n6396 n6394 VDD GND NOR2_X1
xU8979 n8319 n66 n6398 VDD GND NOR2_X1
xU8980 n6456 n6457 n8048 VDD GND NAND2_X1
xU8981 n6461 n6462 n6456 VDD GND NOR2_X1
xU8982 n6458 n6459 n6457 VDD GND NOR2_X1
xU8983 n8320 n75 n6461 VDD GND NOR2_X1
xU8984 n6421 n6422 n8043 VDD GND NAND2_X1
xU8985 n6426 n6427 n6421 VDD GND NOR2_X1
xU8986 n6423 n6424 n6422 VDD GND NOR2_X1
xU8987 n8320 n70 n6426 VDD GND NOR2_X1
xU8988 n6449 n6450 n8047 VDD GND NAND2_X1
xU8989 n6454 n6455 n6449 VDD GND NOR2_X1
xU8990 n6451 n6452 n6450 VDD GND NOR2_X1
xU8991 n8320 n74 n6454 VDD GND NOR2_X1
xU8992 n6288 n6289 n8024 VDD GND NAND2_X1
xU8993 n6293 n6294 n6288 VDD GND NOR2_X1
xU8994 n6290 n6291 n6289 VDD GND NOR2_X1
xU8995 n8318 n51 n6293 VDD GND NOR2_X1
xU8996 n6407 n6408 n8041 VDD GND NAND2_X1
xU8997 n6412 n6413 n6407 VDD GND NOR2_X1
xU8998 n6409 n6410 n6408 VDD GND NOR2_X1
xU8999 n8319 n68 n6412 VDD GND NOR2_X1
xU9000 n6190 n6191 n8010 VDD GND NAND2_X1
xU9001 n6195 n6196 n6190 VDD GND NOR2_X1
xU9002 n6192 n6193 n6191 VDD GND NOR2_X1
xU9003 n8316 n37 n6195 VDD GND NOR2_X1
xU9004 n6414 n6415 n8042 VDD GND NAND2_X1
xU9005 n6419 n6420 n6414 VDD GND NOR2_X1
xU9006 n6416 n6417 n6415 VDD GND NOR2_X1
xU9007 n8319 n69 n6419 VDD GND NOR2_X1
xU9008 n6099 n6100 n7997 VDD GND NAND2_X1
xU9009 n6104 n6105 n6099 VDD GND NOR2_X1
xU9010 n6101 n6102 n6100 VDD GND NOR2_X1
xU9011 n8315 n24 n6104 VDD GND NOR2_X1
xU9012 n6043 n6044 n7989 VDD GND NAND2_X1
xU9013 n6048 n6049 n6043 VDD GND NOR2_X1
xU9014 n6045 n6046 n6044 VDD GND NOR2_X1
xU9015 n8314 n16 n6048 VDD GND NOR2_X1
xU9016 n6036 n6037 n7988 VDD GND NAND2_X1
xU9017 n6041 n6042 n6036 VDD GND NOR2_X1
xU9018 n6038 n6039 n6037 VDD GND NOR2_X1
xU9019 n8314 n15 n6041 VDD GND NOR2_X1
xU9020 n5973 n5974 n7979 VDD GND NAND2_X1
xU9021 n5978 n5979 n5973 VDD GND NOR2_X1
xU9022 n5975 n5976 n5974 VDD GND NOR2_X1
xU9023 n8313 n6 n5978 VDD GND NOR2_X1
xU9024 n6008 n6009 n7984 VDD GND NAND2_X1
xU9025 n6013 n6014 n6008 VDD GND NOR2_X1
xU9026 n6010 n6011 n6009 VDD GND NOR2_X1
xU9027 n8314 n11 n6013 VDD GND NOR2_X1
xU9028 n7394 n7395 n8099 VDD GND NAND2_X1
xU9029 n7422 n7423 n7394 VDD GND NOR2_X1
xU9030 n7396 n7397 n7395 VDD GND NOR2_X1
xU9031 n8325 n126 n7423 VDD GND NOR2_X1
xU9032 n6064 n6065 n7992 VDD GND NAND2_X1
xU9033 n6069 n6070 n6064 VDD GND NOR2_X1
xU9034 n6066 n6067 n6065 VDD GND NOR2_X1
xU9035 n8314 n19 n6069 VDD GND NOR2_X1
xU9036 n5966 n5967 n7978 VDD GND NAND2_X1
xU9037 n5971 n5972 n5966 VDD GND NOR2_X1
xU9038 n5968 n5969 n5967 VDD GND NOR2_X1
xU9039 n8313 n5 n5971 VDD GND NOR2_X1
xU9040 n8329 n6607 n6605 VDD GND NOR2_X1
xU9041 n8329 n6565 n6563 VDD GND NOR2_X1
xU9042 n8329 n6509 n6507 VDD GND NOR2_X1
xU9043 n8329 n6572 n6570 VDD GND NOR2_X1
xU9044 n8329 n6516 n6514 VDD GND NOR2_X1
xU9045 n8329 n6600 n6598 VDD GND NOR2_X1
xU9046 n8329 n6488 n6486 VDD GND NOR2_X1
xU9047 n8329 n6544 n6542 VDD GND NOR2_X1
xU9048 n8329 n6495 n6493 VDD GND NOR2_X1
xU9049 n8329 n6551 n6549 VDD GND NOR2_X1
xU9050 n4569 n488 VDD GND INV_X1
xU9051 n5703 n5699 n5690 VDD GND NAND2_X1
xU9052 n4657 n461 VDD GND INV_X1
xU9053 n3422 n247 VDD GND INV_X1
xU9054 n5609 n5622 n5377 VDD GND NAND2_X1
xU9055 n5987 n5988 n7981 VDD GND NAND2_X1
xU9056 n5992 n5993 n5987 VDD GND NOR2_X1
xU9057 n5989 n5990 n5988 VDD GND NOR2_X1
xU9058 n8313 n8 n5992 VDD GND NOR2_X1
xU9059 n6127 n6128 n8001 VDD GND NAND2_X1
xU9060 n6132 n6133 n6127 VDD GND NOR2_X1
xU9061 n6129 n6130 n6128 VDD GND NOR2_X1
xU9062 n8315 n28 n6132 VDD GND NOR2_X1
xU9063 n5980 n5981 n7980 VDD GND NAND2_X1
xU9064 n5985 n5986 n5980 VDD GND NOR2_X1
xU9065 n5982 n5983 n5981 VDD GND NOR2_X1
xU9066 n8313 n7 n5985 VDD GND NOR2_X1
xU9067 n6022 n6023 n7986 VDD GND NAND2_X1
xU9068 n6027 n6028 n6022 VDD GND NOR2_X1
xU9069 n6024 n6025 n6023 VDD GND NOR2_X1
xU9070 n8314 n13 n6027 VDD GND NOR2_X1
xU9071 n6078 n6079 n7994 VDD GND NAND2_X1
xU9072 n6083 n6084 n6078 VDD GND NOR2_X1
xU9073 n6080 n6081 n6079 VDD GND NOR2_X1
xU9074 n8315 n21 n6083 VDD GND NOR2_X1
xU9075 n6029 n6030 n7987 VDD GND NAND2_X1
xU9076 n6034 n6035 n6029 VDD GND NOR2_X1
xU9077 n6031 n6032 n6030 VDD GND NOR2_X1
xU9078 n8314 n14 n6034 VDD GND NOR2_X1
xU9079 n5936 n5937 n7974 VDD GND NAND2_X1
xU9080 n5942 n5943 n5936 VDD GND NOR2_X1
xU9081 n5938 n5939 n5937 VDD GND NOR2_X1
xU9082 n8319 n1 n5942 VDD GND NOR2_X1
xU9083 n6141 n6142 n8003 VDD GND NAND2_X1
xU9084 n6146 n6147 n6141 VDD GND NOR2_X1
xU9085 n6143 n6144 n6142 VDD GND NOR2_X1
xU9086 n8315 n30 n6146 VDD GND NOR2_X1
xU9087 n6050 n6051 n7990 VDD GND NAND2_X1
xU9088 n6055 n6056 n6050 VDD GND NOR2_X1
xU9089 n6052 n6053 n6051 VDD GND NOR2_X1
xU9090 n8314 n17 n6055 VDD GND NOR2_X1
xU9091 n6071 n6072 n7993 VDD GND NAND2_X1
xU9092 n6076 n6077 n6071 VDD GND NOR2_X1
xU9093 n6073 n6074 n6072 VDD GND NOR2_X1
xU9094 n8314 n20 n6076 VDD GND NOR2_X1
xU9095 n6106 n6107 n7998 VDD GND NAND2_X1
xU9096 n6111 n6112 n6106 VDD GND NOR2_X1
xU9097 n6108 n6109 n6107 VDD GND NOR2_X1
xU9098 n8315 n25 n6111 VDD GND NOR2_X1
xU9099 n6603 n6604 n8069 VDD GND NAND2_X1
xU9100 n6608 n6609 n6603 VDD GND NOR2_X1
xU9101 n6605 n6606 n6604 VDD GND NOR2_X1
xU9102 n8322 n96 n6608 VDD GND NOR2_X1
xU9103 n6351 n6352 n8033 VDD GND NAND2_X1
xU9104 n6356 n6357 n6351 VDD GND NOR2_X1
xU9105 n6353 n6354 n6352 VDD GND NOR2_X1
xU9106 n8318 n60 n6356 VDD GND NOR2_X1
xU9107 n6092 n6093 n7996 VDD GND NAND2_X1
xU9108 n6097 n6098 n6092 VDD GND NOR2_X1
xU9109 n6094 n6095 n6093 VDD GND NOR2_X1
xU9110 n8315 n23 n6097 VDD GND NOR2_X1
xU9111 n6309 n6310 n8027 VDD GND NAND2_X1
xU9112 n6314 n6315 n6309 VDD GND NOR2_X1
xU9113 n6311 n6312 n6310 VDD GND NOR2_X1
xU9114 n8318 n54 n6314 VDD GND NOR2_X1
xU9115 n6358 n6359 n8034 VDD GND NAND2_X1
xU9116 n6363 n6364 n6358 VDD GND NOR2_X1
xU9117 n6360 n6361 n6359 VDD GND NOR2_X1
xU9118 n8319 n61 n6363 VDD GND NOR2_X1
xU9119 n6365 n6366 n8035 VDD GND NAND2_X1
xU9120 n6370 n6371 n6365 VDD GND NOR2_X1
xU9121 n6367 n6368 n6366 VDD GND NOR2_X1
xU9122 n8319 n62 n6370 VDD GND NOR2_X1
xU9123 n6330 n6331 n8030 VDD GND NAND2_X1
xU9124 n6335 n6336 n6330 VDD GND NOR2_X1
xU9125 n6332 n6333 n6331 VDD GND NOR2_X1
xU9126 n8318 n57 n6335 VDD GND NOR2_X1
xU9127 n6554 n6555 n8062 VDD GND NAND2_X1
xU9128 n6559 n6560 n6554 VDD GND NOR2_X1
xU9129 n6556 n6557 n6555 VDD GND NOR2_X1
xU9130 n8321 n89 n6559 VDD GND NOR2_X1
xU9131 n6400 n6401 n8040 VDD GND NAND2_X1
xU9132 n6405 n6406 n6400 VDD GND NOR2_X1
xU9133 n6402 n6403 n6401 VDD GND NOR2_X1
xU9134 n8319 n67 n6405 VDD GND NOR2_X1
xU9135 n6442 n6443 n8046 VDD GND NAND2_X1
xU9136 n6447 n6448 n6442 VDD GND NOR2_X1
xU9137 n6444 n6445 n6443 VDD GND NOR2_X1
xU9138 n8320 n73 n6447 VDD GND NOR2_X1
xU9139 n6463 n6464 n8049 VDD GND NAND2_X1
xU9140 n6468 n6469 n6463 VDD GND NOR2_X1
xU9141 n6465 n6466 n6464 VDD GND NOR2_X1
xU9142 n8320 n76 n6468 VDD GND NOR2_X1
xU9143 n6519 n6520 n8057 VDD GND NAND2_X1
xU9144 n6524 n6525 n6519 VDD GND NOR2_X1
xU9145 n6521 n6522 n6520 VDD GND NOR2_X1
xU9146 n8321 n84 n6524 VDD GND NOR2_X1
xU9147 n6561 n6562 n8063 VDD GND NAND2_X1
xU9148 n6566 n6567 n6561 VDD GND NOR2_X1
xU9149 n6563 n6564 n6562 VDD GND NOR2_X1
xU9150 n8322 n90 n6566 VDD GND NOR2_X1
xU9151 n6498 n6499 n8054 VDD GND NAND2_X1
xU9152 n6503 n6504 n6498 VDD GND NOR2_X1
xU9153 n6500 n6501 n6499 VDD GND NOR2_X1
xU9154 n8321 n81 n6503 VDD GND NOR2_X1
xU9155 n6589 n6590 n8067 VDD GND NAND2_X1
xU9156 n6594 n6595 n6589 VDD GND NOR2_X1
xU9157 n6591 n6592 n6590 VDD GND NOR2_X1
xU9158 n8322 n94 n6594 VDD GND NOR2_X1
xU9159 n6505 n6506 n8055 VDD GND NAND2_X1
xU9160 n6510 n6511 n6505 VDD GND NOR2_X1
xU9161 n6507 n6508 n6506 VDD GND NOR2_X1
xU9162 n8321 n82 n6510 VDD GND NOR2_X1
xU9163 n6568 n6569 n8064 VDD GND NAND2_X1
xU9164 n6573 n6574 n6568 VDD GND NOR2_X1
xU9165 n6570 n6571 n6569 VDD GND NOR2_X1
xU9166 n8322 n91 n6573 VDD GND NOR2_X1
xU9167 n6386 n6387 n8038 VDD GND NAND2_X1
xU9168 n6391 n6392 n6386 VDD GND NOR2_X1
xU9169 n6388 n6389 n6387 VDD GND NOR2_X1
xU9170 n8319 n65 n6391 VDD GND NOR2_X1
xU9171 n6477 n6478 n8051 VDD GND NAND2_X1
xU9172 n6482 n6483 n6477 VDD GND NOR2_X1
xU9173 n6479 n6480 n6478 VDD GND NOR2_X1
xU9174 n8320 n78 n6482 VDD GND NOR2_X1
xU9175 n6526 n6527 n8058 VDD GND NAND2_X1
xU9176 n6531 n6532 n6526 VDD GND NOR2_X1
xU9177 n6528 n6529 n6527 VDD GND NOR2_X1
xU9178 n8321 n85 n6531 VDD GND NOR2_X1
xU9179 n6512 n6513 n8056 VDD GND NAND2_X1
xU9180 n6517 n6518 n6512 VDD GND NOR2_X1
xU9181 n6514 n6515 n6513 VDD GND NOR2_X1
xU9182 n8321 n83 n6517 VDD GND NOR2_X1
xU9183 n6582 n6583 n8066 VDD GND NAND2_X1
xU9184 n6587 n6588 n6582 VDD GND NOR2_X1
xU9185 n6584 n6585 n6583 VDD GND NOR2_X1
xU9186 n8322 n93 n6587 VDD GND NOR2_X1
xU9187 n6470 n6471 n8050 VDD GND NAND2_X1
xU9188 n6475 n6476 n6470 VDD GND NOR2_X1
xU9189 n6472 n6473 n6471 VDD GND NOR2_X1
xU9190 n8320 n77 n6475 VDD GND NOR2_X1
xU9191 n6533 n6534 n8059 VDD GND NAND2_X1
xU9192 n6538 n6539 n6533 VDD GND NOR2_X1
xU9193 n6535 n6536 n6534 VDD GND NOR2_X1
xU9194 n8321 n86 n6538 VDD GND NOR2_X1
xU9195 n6596 n6597 n8068 VDD GND NAND2_X1
xU9196 n6601 n6602 n6596 VDD GND NOR2_X1
xU9197 n6598 n6599 n6597 VDD GND NOR2_X1
xU9198 n8322 n95 n6601 VDD GND NOR2_X1
xU9199 n6428 n6429 n8044 VDD GND NAND2_X1
xU9200 n6433 n6434 n6428 VDD GND NOR2_X1
xU9201 n6430 n6431 n6429 VDD GND NOR2_X1
xU9202 n8320 n71 n6433 VDD GND NOR2_X1
xU9203 n6484 n6485 n8052 VDD GND NAND2_X1
xU9204 n6489 n6490 n6484 VDD GND NOR2_X1
xU9205 n6486 n6487 n6485 VDD GND NOR2_X1
xU9206 n8320 n79 n6489 VDD GND NOR2_X1
xU9207 n6540 n6541 n8060 VDD GND NAND2_X1
xU9208 n6545 n6546 n6540 VDD GND NOR2_X1
xU9209 n6542 n6543 n6541 VDD GND NOR2_X1
xU9210 n8321 n87 n6545 VDD GND NOR2_X1
xU9211 n6575 n6576 n8065 VDD GND NAND2_X1
xU9212 n6580 n6581 n6575 VDD GND NOR2_X1
xU9213 n6577 n6578 n6576 VDD GND NOR2_X1
xU9214 n8322 n92 n6580 VDD GND NOR2_X1
xU9215 n6435 n6436 n8045 VDD GND NAND2_X1
xU9216 n6440 n6441 n6435 VDD GND NOR2_X1
xU9217 n6437 n6438 n6436 VDD GND NOR2_X1
xU9218 n8320 n72 n6440 VDD GND NOR2_X1
xU9219 n6491 n6492 n8053 VDD GND NAND2_X1
xU9220 n6496 n6497 n6491 VDD GND NOR2_X1
xU9221 n6493 n6494 n6492 VDD GND NOR2_X1
xU9222 n8321 n80 n6496 VDD GND NOR2_X1
xU9223 n6547 n6548 n8061 VDD GND NAND2_X1
xU9224 n6552 n6553 n6547 VDD GND NOR2_X1
xU9225 n6549 n6550 n6548 VDD GND NOR2_X1
xU9226 n8321 n88 n6552 VDD GND NOR2_X1
xU9227 n4160 n4309 n3978 VDD GND NAND2_X1
xU9228 n7079 n843 VDD GND INV_X1
xU9229 n2019 n676 VDD GND INV_X1
xU9230 n4686 n464 VDD GND INV_X1
xU9231 n3213 n439 VDD GND INV_X1
xU9232 n3441 n251 VDD GND INV_X1
xU9233 n3384 n3450 n3438 VDD GND NAND2_X1
xU9234 n7502 n877 VDD GND INV_X1
xU9235 n6831 n859 VDD GND INV_X1
xU9236 n359 n5850 n5829 VDD GND NAND2_X1
xU9237 n5489 n359 VDD GND INV_X1
xU9238 n4415 n620 VDD GND INV_X1
xU9239 n4496 n305 VDD GND INV_X1
xU9240 n5403 n5546 n4874 VDD GND NAND2_X1
xU9241 n5428 n5563 n5064 VDD GND NAND2_X1
xU9242 n3228 n3229 n3139 VDD GND NAND2_X1
xU9243 n1948 n1944 n1936 VDD GND NAND2_X1
xU9244 n1927 n2078 n1913 VDD GND NAND2_X1
xU9245 n4388 n4384 n4376 VDD GND NAND2_X1
xU9246 n5866 n5862 n5854 VDD GND NAND2_X1
xU9247 n5633 n5630 n5619 VDD GND NAND2_X1
xU9248 n4556 n4562 n4543 VDD GND NAND2_X1
xU9249 n4623 n457 n4371 VDD GND NAND2_X1
xU9250 n7485 n7483 n7475 VDD GND NAND2_X1
xU9251 n4469 n4466 n4457 VDD GND NAND2_X1
xU9252 n7264 n828 VDD GND INV_X1
xU9253 n2964 n3071 n2791 VDD GND NAND2_X1
xU9254 n2123 n193 VDD GND INV_X1
xU9255 n4438 n624 VDD GND INV_X1
xU9256 n4608 n491 VDD GND INV_X1
xU9257 n5674 n391 VDD GND INV_X1
xU9258 n3281 n596 VDD GND INV_X1
xU9259 n4324 n4368 n3604 VDD GND NAND2_X1
xU9260 n6976 n6977 n8084 VDD GND NAND2_X1
xU9261 n7001 n7002 n6976 VDD GND NOR2_X1
xU9262 n6978 n6979 n6977 VDD GND NOR2_X1
xU9263 n8324 n111 n7002 VDD GND NOR2_X1
xU9264 n6740 n6741 n8076 VDD GND NAND2_X1
xU9265 n6769 n6770 n6740 VDD GND NOR2_X1
xU9266 n6742 n6743 n6741 VDD GND NOR2_X1
xU9267 n8323 n103 n6770 VDD GND NOR2_X1
xU9268 n7224 n7225 n8093 VDD GND NAND2_X1
xU9269 n7316 n7317 n7224 VDD GND NOR2_X1
xU9270 n7226 n7227 n7225 VDD GND NOR2_X1
xU9271 n8325 n120 n7317 VDD GND NOR2_X1
xU9272 n6872 n6873 n8078 VDD GND NAND2_X1
xU9273 n6886 n6887 n6872 VDD GND NOR2_X1
xU9274 n6874 n6875 n6873 VDD GND NOR2_X1
xU9275 n8323 n105 n6887 VDD GND NOR2_X1
xU9276 n6913 n6914 n8081 VDD GND NAND2_X1
xU9277 n6932 n6933 n6913 VDD GND NOR2_X1
xU9278 n6915 n6916 n6914 VDD GND NOR2_X1
xU9279 n8323 n108 n6933 VDD GND NOR2_X1
xU9280 n6611 n6612 n8070 VDD GND NAND2_X1
xU9281 n6626 n6627 n6611 VDD GND NOR2_X1
xU9282 n6613 n6614 n6612 VDD GND NOR2_X1
xU9283 n8322 n97 n6627 VDD GND NOR2_X1
xU9284 n7135 n7136 n8089 VDD GND NAND2_X1
xU9285 n7152 n7153 n7135 VDD GND NOR2_X1
xU9286 n7137 n7138 n7136 VDD GND NOR2_X1
xU9287 n8324 n116 n7153 VDD GND NOR2_X1
xU9288 n6708 n6709 n8075 VDD GND NAND2_X1
xU9289 n6738 n6739 n6708 VDD GND NOR2_X1
xU9290 n6710 n6711 n6709 VDD GND NOR2_X1
xU9291 n8323 n102 n6739 VDD GND NOR2_X1
xU9292 n6946 n6947 n8083 VDD GND NAND2_X1
xU9293 n6974 n6975 n6946 VDD GND NOR2_X1
xU9294 n6948 n6949 n6947 VDD GND NOR2_X1
xU9295 n8324 n110 n6975 VDD GND NOR2_X1
xU9296 n6771 n6772 n8077 VDD GND NAND2_X1
xU9297 n6870 n6871 n6771 VDD GND NOR2_X1
xU9298 n6773 n6774 n6772 VDD GND NOR2_X1
xU9299 n8323 n104 n6871 VDD GND NOR2_X1
xU9300 n7003 n7004 n8085 VDD GND NAND2_X1
xU9301 n7094 n7095 n7003 VDD GND NOR2_X1
xU9302 n7005 n7006 n7004 VDD GND NOR2_X1
xU9303 n8324 n112 n7095 VDD GND NOR2_X1
xU9304 n7195 n7196 n8092 VDD GND NAND2_X1
xU9305 n7222 n7223 n7195 VDD GND NOR2_X1
xU9306 n7197 n7198 n7196 VDD GND NOR2_X1
xU9307 n8324 n119 n7223 VDD GND NOR2_X1
xU9308 n6628 n6629 n8071 VDD GND NAND2_X1
xU9309 n6642 n6643 n6628 VDD GND NOR2_X1
xU9310 n6630 n6631 n6629 VDD GND NOR2_X1
xU9311 n8322 n98 n6643 VDD GND NOR2_X1
xU9312 n7318 n7319 n8094 VDD GND NAND2_X1
xU9313 n7330 n7331 n7318 VDD GND NOR2_X1
xU9314 n7320 n7321 n7319 VDD GND NOR2_X1
xU9315 n8325 n121 n7331 VDD GND NOR2_X1
xU9316 n6900 n6901 n8080 VDD GND NAND2_X1
xU9317 n6911 n6912 n6900 VDD GND NOR2_X1
xU9318 n6902 n6903 n6901 VDD GND NOR2_X1
xU9319 n8323 n107 n6912 VDD GND NOR2_X1
xU9320 n7096 n7097 n8086 VDD GND NAND2_X1
xU9321 n7110 n7111 n7096 VDD GND NOR2_X1
xU9322 n7098 n7099 n7097 VDD GND NOR2_X1
xU9323 n8324 n113 n7111 VDD GND NOR2_X1
xU9324 n7344 n7345 n8096 VDD GND NAND2_X1
xU9325 n7357 n7358 n7344 VDD GND NOR2_X1
xU9326 n7346 n7347 n7345 VDD GND NOR2_X1
xU9327 n8325 n123 n7358 VDD GND NOR2_X1
xU9328 n6663 n6664 n8073 VDD GND NAND2_X1
xU9329 n6690 n6691 n6663 VDD GND NOR2_X1
xU9330 n6665 n6666 n6664 VDD GND NOR2_X1
xU9331 n8323 n100 n6691 VDD GND NOR2_X1
xU9332 n7165 n7166 n8091 VDD GND NAND2_X1
xU9333 n7193 n7194 n7165 VDD GND NOR2_X1
xU9334 n7167 n7168 n7166 VDD GND NOR2_X1
xU9335 n8324 n118 n7194 VDD GND NOR2_X1
xU9336 n7359 n7360 n8097 VDD GND NAND2_X1
xU9337 n7380 n7381 n7359 VDD GND NOR2_X1
xU9338 n7361 n7362 n7360 VDD GND NOR2_X1
xU9339 n8325 n124 n7381 VDD GND NOR2_X1
xU9340 n7445 n7446 n8101 VDD GND NAND2_X1
xU9341 n7542 n7543 n7445 VDD GND NOR2_X1
xU9342 n7447 n7448 n7446 VDD GND NOR2_X1
xU9343 n8325 n128 n7543 VDD GND NOR2_X1
xU9344 n6644 n6645 n8072 VDD GND NAND2_X1
xU9345 n6661 n6662 n6644 VDD GND NOR2_X1
xU9346 n6646 n6647 n6645 VDD GND NOR2_X1
xU9347 n8322 n99 n6662 VDD GND NOR2_X1
xU9348 n7332 n7333 n8095 VDD GND NAND2_X1
xU9349 n7342 n7343 n7332 VDD GND NOR2_X1
xU9350 n7334 n7335 n7333 VDD GND NOR2_X1
xU9351 n8325 n122 n7343 VDD GND NOR2_X1
xU9352 n6888 n6889 n8079 VDD GND NAND2_X1
xU9353 n6898 n6899 n6888 VDD GND NOR2_X1
xU9354 n6890 n6891 n6889 VDD GND NOR2_X1
xU9355 n8323 n106 n6899 VDD GND NOR2_X1
xU9356 n7124 n7125 n8088 VDD GND NAND2_X1
xU9357 n7133 n7134 n7124 VDD GND NOR2_X1
xU9358 n7126 n7127 n7125 VDD GND NOR2_X1
xU9359 n8324 n115 n7134 VDD GND NOR2_X1
xU9360 n7112 n7113 n8087 VDD GND NAND2_X1
xU9361 n7122 n7123 n7112 VDD GND NOR2_X1
xU9362 n7114 n7115 n7113 VDD GND NOR2_X1
xU9363 n8324 n114 n7123 VDD GND NOR2_X1
xU9364 n6692 n6693 n8074 VDD GND NAND2_X1
xU9365 n6706 n6707 n6692 VDD GND NOR2_X1
xU9366 n6694 n6695 n6693 VDD GND NOR2_X1
xU9367 n8323 n101 n6707 VDD GND NOR2_X1
xU9368 n5959 n5960 n7977 VDD GND NAND2_X1
xU9369 n5964 n5965 n5959 VDD GND NOR2_X1
xU9370 n5961 n5962 n5960 VDD GND NOR2_X1
xU9371 n8313 n4 n5964 VDD GND NOR2_X1
xU9372 n5952 n5953 n7976 VDD GND NAND2_X1
xU9373 n5957 n5958 n5952 VDD GND NOR2_X1
xU9374 n5954 n5955 n5953 VDD GND NOR2_X1
xU9375 n8313 n3 n5957 VDD GND NOR2_X1
xU9376 n7154 n7155 n8090 VDD GND NAND2_X1
xU9377 n7163 n7164 n7154 VDD GND NOR2_X1
xU9378 n7156 n7157 n7155 VDD GND NOR2_X1
xU9379 n8324 n117 n7164 VDD GND NOR2_X1
xU9380 n7382 n7383 n8098 VDD GND NAND2_X1
xU9381 n7392 n7393 n7382 VDD GND NOR2_X1
xU9382 n7384 n7385 n7383 VDD GND NOR2_X1
xU9383 n8325 n125 n7393 VDD GND NOR2_X1
xU9384 n6934 n6935 n8082 VDD GND NAND2_X1
xU9385 n6944 n6945 n6934 VDD GND NOR2_X1
xU9386 n6936 n6937 n6935 VDD GND NOR2_X1
xU9387 n8323 n109 n6945 VDD GND NOR2_X1
xU9388 n6211 n6212 n8013 VDD GND NAND2_X1
xU9389 n6216 n6217 n6211 VDD GND NOR2_X1
xU9390 n6213 n6214 n6212 VDD GND NOR2_X1
xU9391 n8316 n40 n6216 VDD GND NOR2_X1
xU9392 n6204 n6205 n8012 VDD GND NAND2_X1
xU9393 n6209 n6210 n6204 VDD GND NOR2_X1
xU9394 n6206 n6207 n6205 VDD GND NOR2_X1
xU9395 n8316 n39 n6209 VDD GND NOR2_X1
xU9396 n6085 n6086 n7995 VDD GND NAND2_X1
xU9397 n6090 n6091 n6085 VDD GND NOR2_X1
xU9398 n6087 n6088 n6086 VDD GND NOR2_X1
xU9399 n8315 n22 n6090 VDD GND NOR2_X1
xU9400 n6246 n6247 n8018 VDD GND NAND2_X1
xU9401 n6251 n6252 n6246 VDD GND NOR2_X1
xU9402 n6248 n6249 n6247 VDD GND NOR2_X1
xU9403 n8317 n45 n6251 VDD GND NOR2_X1
xU9404 n6302 n6303 n8026 VDD GND NAND2_X1
xU9405 n6307 n6308 n6302 VDD GND NOR2_X1
xU9406 n6304 n6305 n6303 VDD GND NOR2_X1
xU9407 n8318 n53 n6307 VDD GND NOR2_X1
xU9408 n6253 n6254 n8019 VDD GND NAND2_X1
xU9409 n6258 n6259 n6253 VDD GND NOR2_X1
xU9410 n6255 n6256 n6254 VDD GND NOR2_X1
xU9411 n8317 n46 n6258 VDD GND NOR2_X1
xU9412 n6162 n6163 n8006 VDD GND NAND2_X1
xU9413 n6167 n6168 n6162 VDD GND NOR2_X1
xU9414 n6164 n6165 n6163 VDD GND NOR2_X1
xU9415 n8316 n33 n6167 VDD GND NOR2_X1
xU9416 n6274 n6275 n8022 VDD GND NAND2_X1
xU9417 n6279 n6280 n6274 VDD GND NOR2_X1
xU9418 n6276 n6277 n6275 VDD GND NOR2_X1
xU9419 n8317 n49 n6279 VDD GND NOR2_X1
xU9420 n6295 n6296 n8025 VDD GND NAND2_X1
xU9421 n6300 n6301 n6295 VDD GND NOR2_X1
xU9422 n6297 n6298 n6296 VDD GND NOR2_X1
xU9423 n8318 n52 n6300 VDD GND NOR2_X1
xU9424 n5994 n5995 n7982 VDD GND NAND2_X1
xU9425 n5999 n6000 n5994 VDD GND NOR2_X1
xU9426 n5996 n5997 n5995 VDD GND NOR2_X1
xU9427 n8313 n9 n5999 VDD GND NOR2_X1
xU9428 n6218 n6219 n8014 VDD GND NAND2_X1
xU9429 n6223 n6224 n6218 VDD GND NOR2_X1
xU9430 n6220 n6221 n6219 VDD GND NOR2_X1
xU9431 n8317 n41 n6223 VDD GND NOR2_X1
xU9432 n6176 n6177 n8008 VDD GND NAND2_X1
xU9433 n6181 n6182 n6176 VDD GND NOR2_X1
xU9434 n6178 n6179 n6177 VDD GND NOR2_X1
xU9435 n8316 n35 n6181 VDD GND NOR2_X1
xU9436 n6015 n6016 n7985 VDD GND NAND2_X1
xU9437 n6020 n6021 n6015 VDD GND NOR2_X1
xU9438 n6017 n6018 n6016 VDD GND NOR2_X1
xU9439 n8314 n12 n6020 VDD GND NOR2_X1
xU9440 n6239 n6240 n8017 VDD GND NAND2_X1
xU9441 n6244 n6245 n6239 VDD GND NOR2_X1
xU9442 n6241 n6242 n6240 VDD GND NOR2_X1
xU9443 n8317 n44 n6244 VDD GND NOR2_X1
xU9444 n7424 n7425 n8100 VDD GND NAND2_X1
xU9445 n7443 n7444 n7424 VDD GND NOR2_X1
xU9446 n7426 n7427 n7425 VDD GND NOR2_X1
xU9447 n8325 n127 n7444 VDD GND NOR2_X1
xU9448 n5415 n5573 n5252 VDD GND NAND2_X1
xU9449 n7018 n7019 n6885 VDD GND NAND2_X1
xU9450 n3019 n3020 n2959 VDD GND NAND2_X1
xU9451 n3141 n3156 n2931 VDD GND NAND2_X1
xU9452 n2953 n3103 n2596 VDD GND NAND2_X1
xU9453 n3157 n3200 n3174 VDD GND NAND2_X1
xU9454 n5565 n5566 n5259 VDD GND NAND2_X1
xU9455 n5549 n5550 n5062 VDD GND NAND2_X1
xU9456 n7236 n7237 n7105 VDD GND NAND2_X1
xU9457 n3307 n3089 n2864 VDD GND NAND2_X1
xU9458 n2935 n3075 n2390 VDD GND NAND2_X1
xU9459 n4538 n4636 n4105 VDD GND NAND2_X1
xU9460 n1832 n1833 n1349 VDD GND NAND2_X1
xU9461 n6990 n6991 n6972 VDD GND NAND2_X1
xU9462 n1883 n1916 n1854 VDD GND NAND2_X1
xU9463 n7418 n7419 n7329 VDD GND NAND2_X1
xU9464 n7439 n7464 n7355 VDD GND NAND2_X1
xU9465 n6756 n6795 n6659 VDD GND NAND2_X1
xU9466 n5899 n648 VDD GND INV_X1
xU9467 n6970 n6971 n6881 VDD GND NAND2_X1
xU9468 n2043 n672 VDD GND INV_X1
xU9469 n5383 n5536 n5261 VDD GND NAND2_X1
xU9470 n6792 n6793 n6660 VDD GND NAND2_X1
xU9471 n6736 n6737 n6622 VDD GND NAND2_X1
xU9472 n5692 n5697 n5358 VDD GND NAND2_X1
xU9473 n4538 n4539 n4192 VDD GND NAND2_X1
xU9474 n3021 n3022 n2860 VDD GND NAND2_X1
xU9475 n4315 n4393 n4135 VDD GND NAND2_X1
xU9476 n1832 n2156 n1647 VDD GND NAND2_X1
xU9477 n5549 n5871 n5354 VDD GND NAND2_X1
xU9478 n1883 n1884 n1635 VDD GND NAND2_X1
xU9479 n2135 n2145 n1646 VDD GND NAND2_X1
xU9480 n4455 n4463 n4129 VDD GND NAND2_X1
xU9481 n3121 n3137 n2882 VDD GND NAND2_X1
xU9482 n4357 n4541 n4122 VDD GND NAND2_X1
xU9483 n4272 n4273 n4099 VDD GND NAND2_X1
xU9484 n1933 n1942 n1641 VDD GND NAND2_X1
xU9485 n4374 n4382 n4134 VDD GND NAND2_X1
xU9486 n1878 n1911 n1634 VDD GND NAND2_X1
xU9487 n7461 n7462 n7356 VDD GND NAND2_X1
xU9488 n3379 n3399 n2888 VDD GND NAND2_X1
xU9489 n7015 n7016 n6883 VDD GND NAND2_X1
xU9490 n5565 n5708 n5359 VDD GND NAND2_X1
xU9491 n3079 n3148 n2893 VDD GND NAND2_X1
xU9492 n3307 n3316 n2966 VDD GND NAND2_X1
xU9493 n6990 n7020 n6910 VDD GND NAND2_X1
xU9494 n1894 n1895 n1702 VDD GND NAND2_X1
xU9495 n7244 n7245 n7109 VDD GND NAND2_X1
xU9496 n1686 n1857 n1520 VDD GND NAND2_X1
xU9497 n5893 n5873 n5870 VDD GND NAND2_X1
xU9498 n5906 n642 VDD GND INV_X1
xU9499 n3094 n3385 n2889 VDD GND NAND2_X1
xU9500 n4329 n4474 n4130 VDD GND NAND2_X1
xU9501 n4360 n4361 n4123 VDD GND NAND2_X1
xU9502 n4579 n4561 n4559 VDD GND NAND2_X1
xU9503 n7492 n881 VDD GND INV_X1
xU9504 n2049 n675 VDD GND INV_X1
xU9505 n1844 n1953 n1642 VDD GND NAND2_X1
xU9506 n6827 n862 VDD GND INV_X1
xU9507 n3185 n438 VDD GND INV_X1
xU9508 n4408 n623 VDD GND INV_X1
xU9509 n6790 n6791 n6689 VDD GND NAND2_X1
xU9510 n4204 n4321 n4035 VDD GND NAND2_X1
xU9511 n4186 n4320 n4020 VDD GND NAND2_X1
xU9512 n1939 n2005 n1985 VDD GND NAND2_X1
xU9513 n5780 n5781 n5418 VDD GND NAND2_X1
xU9514 n5600 n5601 n5347 VDD GND NAND2_X1
xU9515 n1803 n1804 n1617 VDD GND NAND2_X1
xU9516 n4489 n308 VDD GND INV_X1
xU9517 n1715 n1830 n1152 VDD GND AND2_X1
xU9518 n7207 n7208 n7205 VDD GND NAND2_X1
xU9519 n7374 n7442 n7415 VDD GND NAND2_X1
xU9520 n6964 n7023 n6943 VDD GND NAND2_X1
xU9521 n7412 n7471 n7391 VDD GND NAND2_X1
xU9522 n3407 n3401 n3398 VDD GND NAND2_X1
xU9523 n3410 n250 VDD GND INV_X1
xU9524 n5652 n5624 n5638 VDD GND NAND2_X1
xU9525 n5663 n385 VDD GND INV_X1
xU9526 n6687 n6762 n6735 VDD GND NAND2_X1
xU9527 n4286 n4537 n3951 VDD GND NAND2_X1
xU9528 n3436 n3394 n3406 VDD GND NAND2_X1
xU9529 n3036 n3147 n2939 VDD GND NAND2_X1
xU9530 n4267 n4386 n4190 VDD GND NAND2_X1
xU9531 n6726 n6783 n6705 VDD GND NAND2_X1
xU9532 n3045 n3350 n3364 VDD GND NAND2_X1
xU9533 n6930 n6995 n6967 VDD GND NAND2_X1
xU9534 n1780 n2149 n1718 VDD GND NAND2_X1
xU9535 n5544 n380 VDD GND INV_X1
xU9536 n1764 n1882 n1674 VDD GND NAND2_X1
xU9537 n3010 n3125 n2922 VDD GND NAND2_X1
xU9538 n3262 n3244 n3235 VDD GND NAND2_X1
xU9539 n2095 n2077 n1930 VDD GND NAND2_X1
xU9540 n1978 n1955 n1952 VDD GND NAND2_X1
xU9541 n1989 n410 VDD GND INV_X1
xU9542 n7056 n7029 n7042 VDD GND NAND2_X1
xU9543 n6837 n6803 n6813 VDD GND NAND2_X1
xU9544 n6847 n856 VDD GND INV_X1
xU9545 n6814 n6815 n6807 VDD GND NAND2_X1
xU9546 n4325 n481 VDD GND INV_X1
xU9547 n3390 n237 VDD GND INV_X1
xU9548 n5830 n5791 n5787 VDD GND NAND2_X1
xU9549 n1775 n1892 n1468 VDD GND NAND2_X1
xU9550 n7043 n7039 n7033 VDD GND NAND2_X1
xU9551 n3247 n3248 n3234 VDD GND NAND2_X1
xU9552 n2105 n1926 n2082 VDD GND NAND2_X1
xU9553 n5909 n5863 n5881 VDD GND NAND2_X1
xU9554 n587 n3135 n2914 VDD GND NAND2_X1
xU9555 n3136 n587 VDD GND INV_X1
xU9556 n7508 n873 n7487 VDD GND NAND2_X1
xU9557 n2046 n666 VDD GND INV_X1
xU9558 n2180 n534 n2155 VDD GND NAND2_X1
xU9559 n4405 n614 VDD GND INV_X1
xU9560 n7509 n873 VDD GND INV_X1
xU9561 n3046 n3047 n2961 VDD GND NAND2_X1
xU9562 n615 n4396 n4392 VDD GND NAND2_X1
xU9563 n4425 n615 VDD GND INV_X1
xU9564 n2151 n2147 n2139 VDD GND OR2_X1
xU9565 n5510 n5511 n5400 VDD GND NAND2_X1
xU9566 n5689 n5694 n5422 VDD GND AND2_X1
xU9567 n1963 n1957 n1951 VDD GND NAND2_X1
xU9568 n4485 n4476 n4472 VDD GND NAND2_X1
xU9569 n7488 n7482 n7479 VDD GND NAND2_X1
xU9570 n4647 n4638 n4634 VDD GND NAND2_X1
xU9571 n7298 n821 n7257 VDD GND NAND2_X1
xU9572 n5811 n358 VDD GND INV_X1
xU9573 n5853 n5857 n5396 VDD GND AND2_X1
xU9574 n2137 n2142 n1709 VDD GND AND2_X1
xU9575 n1935 n1939 n1690 VDD GND AND2_X1
xU9576 n4456 n4460 n4198 VDD GND AND2_X1
xU9577 n4270 n4271 n4170 VDD GND AND2_X1
xU9578 n4318 n4317 n4181 VDD GND AND2_X1
xU9579 n1890 n1891 n1681 VDD GND AND2_X1
xU9580 n3135 n3290 n3271 VDD GND AND2_X1
xU9581 n5694 n5766 n5757 VDD GND AND2_X1
xU9582 n6791 n6863 n6843 VDD GND AND2_X1
xU9583 n7460 n7539 n7516 VDD GND AND2_X1
xU9584 n7019 n7081 n7064 VDD GND AND2_X1
xU9585 n3156 n3221 n3203 VDD GND AND2_X1
xU9586 n5622 n5684 n5675 VDD GND AND2_X1
xU9587 n7237 n7312 n7276 VDD GND AND2_X1
xU9588 n4379 n4447 n4427 VDD GND AND2_X1
xU9589 n4271 n4693 n4670 VDD GND AND2_X1
xU9590 n4460 n4530 n4510 VDD GND AND2_X1
xU9591 n4540 n4616 n4586 VDD GND AND2_X1
xU9592 n3393 n3455 n3445 VDD GND AND2_X1
xU9593 n1910 n2127 n2118 VDD GND AND2_X1
xU9594 n2142 n2210 n2187 VDD GND AND2_X1
xU9595 n1802 n2067 n2034 VDD GND AND2_X1
xU9596 n5571 n5569 n5423 VDD GND AND2_X1
xU9597 n3380 n3393 n2947 VDD GND AND2_X1
xU9598 n1801 n1802 n1680 VDD GND AND2_X1
xU9599 n3342 n3306 n3326 VDD GND AND2_X1
xU9600 n3020 n3376 n3365 VDD GND AND2_X1
xU9601 n5857 n5928 n5908 VDD GND AND2_X1
xU9602 n5600 n5610 n5542 VDD GND AND2_X1
xU9603 n4360 n4545 n4339 VDD GND AND2_X1
xU9604 n1844 n1845 n1545 VDD GND AND2_X1
xU9605 n3126 n3236 n3101 VDD GND AND2_X1
xU9606 n479 n4540 n4154 VDD GND AND2_X1
xU9607 n613 n4379 n4180 VDD GND AND2_X1
xU9608 n183 n1910 n1665 VDD GND AND2_X1
xU9609 n3352 n3323 n3315 VDD GND AND2_X1
xU9610 n5852 n5860 n5353 VDD GND AND2_X1
xU9611 n5593 n5629 n5346 VDD GND AND2_X1
xU9612 n3145 n3162 n2892 VDD GND AND2_X1
xU9613 n5490 n5491 n5330 VDD GND AND2_X1
xU9614 n3126 n3127 n2883 VDD GND AND2_X1
xU9615 n5727 n509 VDD GND INV_X1
xU9616 n5720 n5710 n5706 VDD GND AND2_X1
xU9617 n7150 n7216 n7178 VDD GND AND2_X1
xU9618 n4663 n4640 n4635 VDD GND OR2_X1
xU9619 n4502 n4477 n4473 VDD GND OR2_X1
xU9620 n3267 n592 VDD GND INV_X1
xU9621 n2101 n189 VDD GND INV_X1
xU9622 n5397 n639 VDD GND INV_X1
xU9623 n5402 n5403 n5401 VDD GND NAND2_X1
xU9624 n2024 n2025 n1908 VDD GND OR2_X1
xU9625 n6558 n8338 n6556 VDD GND AND2_X1
xU9626 n6404 n8336 n6402 VDD GND AND2_X1
xU9627 n6446 n8337 n6444 VDD GND AND2_X1
xU9628 n6467 n8337 n6465 VDD GND AND2_X1
xU9629 n6523 n8337 n6521 VDD GND AND2_X1
xU9630 n6502 n8337 n6500 VDD GND AND2_X1
xU9631 n6593 n8338 n6591 VDD GND AND2_X1
xU9632 n6390 n8336 n6388 VDD GND AND2_X1
xU9633 n6481 n8337 n6479 VDD GND AND2_X1
xU9634 n6530 n8337 n6528 VDD GND AND2_X1
xU9635 n6586 n8338 n6584 VDD GND AND2_X1
xU9636 n6474 n8337 n6472 VDD GND AND2_X1
xU9637 n6537 n8337 n6535 VDD GND AND2_X1
xU9638 n6432 n8336 n6430 VDD GND AND2_X1
xU9639 n6579 n8338 n6577 VDD GND AND2_X1
xU9640 n6439 n8337 n6437 VDD GND AND2_X1
xU9641 n1914 n184 VDD GND INV_X1
xU9642 n3270 n590 VDD GND INV_X1
xU9643 n2117 n186 VDD GND INV_X1
xU9644 n5911 n646 VDD GND INV_X1
xU9645 n2211 n536 VDD GND INV_X1
xU9646 n6313 n8336 n6311 VDD GND AND2_X1
xU9647 n6222 n8335 n6220 VDD GND AND2_X1
xU9648 n6180 n8335 n6178 VDD GND AND2_X1
xU9649 n6243 n8335 n6241 VDD GND AND2_X1
xU9650 n5956 n8337 n5954 VDD GND AND2_X1
xU9651 n5998 n8334 n5996 VDD GND AND2_X1
xU9652 n6215 n8335 n6213 VDD GND AND2_X1
xU9653 n6355 n8336 n6353 VDD GND AND2_X1
xU9654 n6208 n8335 n6206 VDD GND AND2_X1
xU9655 n6250 n8335 n6248 VDD GND AND2_X1
xU9656 n6362 n8336 n6360 VDD GND AND2_X1
xU9657 n6306 n8336 n6304 VDD GND AND2_X1
xU9658 n6257 n8335 n6255 VDD GND AND2_X1
xU9659 n6166 n8335 n6164 VDD GND AND2_X1
xU9660 n6369 n8336 n6367 VDD GND AND2_X1
xU9661 n6278 n8335 n6276 VDD GND AND2_X1
xU9662 n6299 n8336 n6297 VDD GND AND2_X1
xU9663 n6334 n8336 n6332 VDD GND AND2_X1
xU9664 n8340 n6096 n6094 VDD GND AND2_X1
xU9665 n7452 n131 n7546 VDD GND NOR2_X1
xU9666 n7570 n131 VDD GND INV_X1
xU9667 n8326 n6061 n6059 VDD GND NOR2_X1
xU9668 n8326 n6005 n6003 VDD GND NOR2_X1
xU9669 n8326 n5949 n5947 VDD GND NOR2_X1
xU9670 n8326 n6117 n6115 VDD GND NOR2_X1
xU9671 n6057 n6058 n7991 VDD GND NAND2_X1
xU9672 n6062 n6063 n6057 VDD GND NOR2_X1
xU9673 n6059 n6060 n6058 VDD GND NOR2_X1
xU9674 n8314 n18 n6062 VDD GND NOR2_X1
xU9675 n6001 n6002 n7983 VDD GND NAND2_X1
xU9676 n6006 n6007 n6001 VDD GND NOR2_X1
xU9677 n6003 n6004 n6002 VDD GND NOR2_X1
xU9678 n8313 n10 n6006 VDD GND NOR2_X1
xU9679 n5945 n5946 n7975 VDD GND NAND2_X1
xU9680 n5950 n5951 n5945 VDD GND NOR2_X1
xU9681 n5947 n5948 n5946 VDD GND NOR2_X1
xU9682 n8313 n2 n5950 VDD GND NOR2_X1
xU9683 n6113 n6114 n7999 VDD GND NAND2_X1
xU9684 n6118 n6119 n6113 VDD GND NOR2_X1
xU9685 n6115 n6116 n6114 VDD GND NOR2_X1
xU9686 n8315 n26 n6118 VDD GND NOR2_X1
xU9687 n6680 n810 VDD GND INV_X1
xU9688 n6641 n811 VDD GND INV_X1
xU9689 n6704 n812 VDD GND INV_X1
xU9690 n6680 n6656 n6765 VDD GND AND2_X1
xU9691 n5935 n8357 n1009 VDD GND NAND2_X1
xU9692 n8362 n7451 n6610 VDD GND NOR2_X1
xU9693 n135 n7452 n7451 VDD GND NOR2_X1
xU9694 n5944 n8310 VDD GND BUF_X1
xU9695 n5944 n8311 VDD GND BUF_X1
xU9696 n7579 n8256 VDD GND BUF_X1
xU9697 n7579 n8255 VDD GND BUF_X1
xU9698 n989 n8399 VDD GND BUF_X1
xU9699 n989 n8400 VDD GND BUF_X1
xU9700 n989 n8401 VDD GND BUF_X1
xU9701 n5944 n8312 VDD GND BUF_X1
xU9702 n7579 n8257 VDD GND BUF_X1
xU9703 n7578 n8271 VDD GND BUF_X1
xU9704 n7452 n8258 n7578 VDD GND NOR2_X1
xU9705 n7839 n130 VDD GND INV_X1
xU9706 n7452 n136 VDD GND INV_X1
xU9707 n7455 n133 VDD GND INV_X1
xU9708 n6640 \AES_Comp_ENCa/Rrg_6 n6639 VDD GND NAND2_X1
xU9709 n6703 n810 n6701 VDD GND NOR2_X1
xU9710 n5837 n5573 n5836 VDD GND NAND2_X1
xU9711 n1714 n1715 n1713 VDD GND NAND2_X1
xU9712 n1895 n2051 n2036 VDD GND NAND2_X1
xU9713 n4326 n4674 n4651 VDD GND NAND2_X1
xU9714 n3103 n3448 n3412 VDD GND NAND2_X1
xU9715 n2961 n8252 n8251 VDD GND XOR2_X1
xU9716 n2963 n560 n8252 VDD GND OR2_X1
xU9717 n1695 n1696 n1694 VDD GND NAND2_X1
xU9718 n1685 n1686 n1684 VDD GND NAND2_X1
xU9719 n4203 n4204 n4202 VDD GND NAND2_X1
xU9720 n5427 n5428 n5426 VDD GND NAND2_X1
xU9721 n5382 n5383 n5381 VDD GND NAND2_X1
xU9722 n2952 n2953 n2951 VDD GND NAND2_X1
xU9723 n1670 n1671 n1669 VDD GND NAND2_X1
xU9724 n4159 n4160 n4158 VDD GND NAND2_X1
xU9725 n4185 n4186 n4184 VDD GND NAND2_X1
xU9726 n872 n7372 n7370 VDD GND NOR2_X1
xU9727 n7374 n872 VDD GND INV_X1
xU9728 n810 \AES_Comp_ENCa/Rrg_0 n6781 VDD GND NOR2_X1
xU9729 n6656 n6657 n6655 VDD GND NAND2_X1
xU9730 \AES_Comp_ENCa/Rrg_5 n811 n6657 VDD GND NAND2_X1
xU9731 n6656 n6730 n6728 VDD GND NAND2_X1
xU9732 n6731 \AES_Comp_ENCa/Rrg_2 n6730 VDD GND NAND2_X1
xU9733 \AES_Comp_ENCa/Rrg_1 \AES_Comp_ENCa/Rrg_0 n6731 VDD GND NOR2_X1
xU9734 n6678 n6679 n6677 VDD GND NOR2_X1
xU9735 n815 n6681 n6678 VDD GND NOR2_X1
xU9736 n6656 n6680 n6679 VDD GND NAND2_X1
xU9737 n8326 n7400 n7396 VDD GND NOR2_X1
xU9738 n6593 n826 n7400 VDD GND NAND2_X1
xU9739 Dout_E_62 n4684 n4652 VDD GND AND2_X1
xU9740 n362 n5488 n5328 VDD GND NOR2_X1
xU9741 n593 n3136 n3128 VDD GND NOR2_X1
xU9742 n618 n4375 n4314 VDD GND NOR2_X1
xU9743 n3071 n3360 n3353 VDD GND AND2_X1
xU9744 n485 n4544 n4358 VDD GND NOR2_X1
xU9745 n190 n1915 n1880 VDD GND NOR2_X1
xU9746 n3207 n3075 n3187 VDD GND AND2_X1
xU9747 n5560 n5561 n4719 VDD GND NAND2_X1
xU9748 n1846 n1847 n1244 VDD GND NAND2_X1
xU9749 n5567 n5568 n4962 VDD GND NAND2_X1
xU9750 n4330 n4331 n3531 VDD GND NAND2_X1
xU9751 n5551 n5552 n4770 VDD GND NAND2_X1
xU9752 n4627 n4624 n4104 VDD GND NAND2_X1
xU9753 n1834 n1835 n1050 VDD GND NAND2_X1
xU9754 n5693 n5744 n5727 VDD GND NAND2_X1
xU9755 n1920 n185 n1437 VDD GND NAND2_X1
xU9756 n4316 n611 n3725 VDD GND NAND2_X1
xU9757 n1899 n1896 n1613 VDD GND NAND2_X1
xU9758 n5604 n5605 n4873 VDD GND NAND2_X1
xU9759 n4537 n4681 n4665 VDD GND NAND2_X1
xU9760 n3125 n3283 n3264 VDD GND NAND2_X1
xU9761 n1882 n2102 n2089 VDD GND NAND2_X1
xU9762 n7471 n7529 n7511 VDD GND NAND2_X1
xU9763 n4321 n4514 n4490 VDD GND NAND2_X1
xU9764 n7023 n7072 n7058 VDD GND NAND2_X1
xU9765 n6783 n6856 n6839 VDD GND NAND2_X1
xU9766 n1946 n1998 n1980 VDD GND NAND2_X1
xU9767 n7442 n7520 n7493 VDD GND NAND2_X1
xU9768 n6762 n6848 n6829 VDD GND NAND2_X1
xU9769 \AES_Comp_ENCa/KrgX_1 n5532 n5526 VDD GND NOR2_X1
xU9770 n5533 n5534 n5532 VDD GND NOR2_X1
xU9771 n8433 n379 n5534 VDD GND NOR2_X1
xU9772 n8398 n5531 n5533 VDD GND NOR2_X1
xU9773 n5864 n5920 n5907 VDD GND NAND2_X1
xU9774 n6980 n857 n6979 VDD GND NOR2_X1
xU9775 n6981 n8298 n6980 VDD GND NOR2_X1
xU9776 n6488 n8339 n6981 VDD GND AND2_X1
xU9777 \AES_Comp_ENCa/KrgX_25 n7459 n7414 VDD GND NAND2_X1
xU9778 n3095 n3096 n2490 VDD GND AND2_X1
xU9779 n6917 n864 n6916 VDD GND NOR2_X1
xU9780 n6918 n8296 n6917 VDD GND NOR2_X1
xU9781 n8328 n6467 n6918 VDD GND NOR2_X1
xU9782 n7322 n832 n7321 VDD GND NOR2_X1
xU9783 n7323 n8303 n7322 VDD GND NOR2_X1
xU9784 n8331 n6558 n7323 VDD GND NOR2_X1
xU9785 n8331 n7324 n7320 VDD GND NOR2_X1
xU9786 n6558 n832 n7324 VDD GND NAND2_X1
xU9787 n6648 n882 n6647 VDD GND NOR2_X1
xU9788 n6649 n8292 n6648 VDD GND NOR2_X1
xU9789 n8329 n6404 n6649 VDD GND NOR2_X1
xU9790 n8330 n6650 n6646 VDD GND NOR2_X1
xU9791 n6404 n882 n6650 VDD GND NAND2_X1
xU9792 n6876 n867 n6875 VDD GND NOR2_X1
xU9793 n6877 n8295 n6876 VDD GND NOR2_X1
xU9794 n8330 n6446 n6877 VDD GND NOR2_X1
xU9795 n8330 n6878 n6874 VDD GND NOR2_X1
xU9796 n6446 n867 n6878 VDD GND NAND2_X1
xU9797 n8330 n6919 n6915 VDD GND NOR2_X1
xU9798 n6467 n864 n6919 VDD GND NAND2_X1
xU9799 n7139 n844 n7138 VDD GND NOR2_X1
xU9800 n7140 n8300 n7139 VDD GND NOR2_X1
xU9801 n8331 n6523 n7140 VDD GND NOR2_X1
xU9802 n7100 n847 n7099 VDD GND NOR2_X1
xU9803 n7101 n8299 n7100 VDD GND NOR2_X1
xU9804 n8330 n6502 n7101 VDD GND NOR2_X1
xU9805 n8331 n7102 n7098 VDD GND NOR2_X1
xU9806 n6502 n847 n7102 VDD GND NAND2_X1
xU9807 n6615 n884 n6614 VDD GND NOR2_X1
xU9808 n6616 n8291 n6615 VDD GND NOR2_X1
xU9809 n8329 n6390 n6616 VDD GND NOR2_X1
xU9810 n8329 n6617 n6613 VDD GND NOR2_X1
xU9811 n6390 n884 n6617 VDD GND NAND2_X1
xU9812 n6950 n860 n6949 VDD GND NOR2_X1
xU9813 n6951 n8297 n6950 VDD GND NOR2_X1
xU9814 n8330 n6481 n6951 VDD GND NOR2_X1
xU9815 n8330 n6952 n6948 VDD GND NOR2_X1
xU9816 n6481 n860 n6952 VDD GND NAND2_X1
xU9817 n7158 n842 n7157 VDD GND NOR2_X1
xU9818 n7159 n8301 n7158 VDD GND NOR2_X1
xU9819 n8331 n6530 n7159 VDD GND NOR2_X1
xU9820 n8331 n7160 n7156 VDD GND NOR2_X1
xU9821 n6530 n842 n7160 VDD GND NAND2_X1
xU9822 n7386 n827 n7385 VDD GND NOR2_X1
xU9823 n7387 n8305 n7386 VDD GND NOR2_X1
xU9824 n8331 n6586 n7387 VDD GND NOR2_X1
xU9825 n6938 n861 n6937 VDD GND NOR2_X1
xU9826 n6939 n8297 n6938 VDD GND NOR2_X1
xU9827 n8330 n6474 n6939 VDD GND NOR2_X1
xU9828 n7169 n841 n7168 VDD GND NOR2_X1
xU9829 n7170 n8301 n7169 VDD GND NOR2_X1
xU9830 n8331 n6537 n7170 VDD GND NOR2_X1
xU9831 n8331 n7171 n7167 VDD GND NOR2_X1
xU9832 n6537 n841 n7171 VDD GND NAND2_X1
xU9833 n6744 n876 n6743 VDD GND NOR2_X1
xU9834 n6745 n8294 n6744 VDD GND NOR2_X1
xU9835 n8330 n6432 n6745 VDD GND NOR2_X1
xU9836 n8330 n6746 n6742 VDD GND NOR2_X1
xU9837 n6432 n876 n6746 VDD GND NAND2_X1
xU9838 n7363 n829 n7362 VDD GND NOR2_X1
xU9839 n7364 n8304 n7363 VDD GND NOR2_X1
xU9840 n8331 n6579 n7364 VDD GND NOR2_X1
xU9841 n8331 n7365 n7361 VDD GND NOR2_X1
xU9842 n6579 n829 n7365 VDD GND NAND2_X1
xU9843 n6775 n875 n6774 VDD GND NOR2_X1
xU9844 n6776 n8294 n6775 VDD GND NOR2_X1
xU9845 n8330 n6439 n6776 VDD GND NOR2_X1
xU9846 n8330 n6777 n6773 VDD GND NOR2_X1
xU9847 n6439 n875 n6777 VDD GND NAND2_X1
xU9848 n6712 n878 n6711 VDD GND NOR2_X1
xU9849 n6713 n8293 n6712 VDD GND NOR2_X1
xU9850 n6425 n8338 n6713 VDD GND AND2_X1
xU9851 n7007 n854 n7006 VDD GND NOR2_X1
xU9852 n7008 n8298 n7007 VDD GND NOR2_X1
xU9853 n6495 n8339 n7008 VDD GND AND2_X1
xU9854 n7199 n840 n7198 VDD GND NOR2_X1
xU9855 n7200 n8302 n7199 VDD GND NOR2_X1
xU9856 n6544 n8339 n7200 VDD GND AND2_X1
xU9857 n3080 n3081 n2281 VDD GND AND2_X1
xU9858 n6600 n7430 n7426 VDD GND NOR2_X1
xU9859 n8332 n825 n7430 VDD GND NAND2_X1
xU9860 n6565 n7338 n7334 VDD GND NOR2_X1
xU9861 n8332 n831 n7338 VDD GND NAND2_X1
xU9862 n6397 n6634 n6630 VDD GND NOR2_X1
xU9863 n8334 n883 n6634 VDD GND NAND2_X1
xU9864 n6460 n6906 n6902 VDD GND NOR2_X1
xU9865 n8333 n865 n6906 VDD GND NAND2_X1
xU9866 n6425 n6714 n6710 VDD GND NOR2_X1
xU9867 n8334 n878 n6714 VDD GND NAND2_X1
xU9868 n6453 n6894 n6890 VDD GND NOR2_X1
xU9869 n8334 n866 n6894 VDD GND NAND2_X1
xU9870 n6509 n7118 n7114 VDD GND NOR2_X1
xU9871 n8332 n846 n7118 VDD GND NAND2_X1
xU9872 n6572 n7350 n7346 VDD GND NOR2_X1
xU9873 n8332 n830 n7350 VDD GND NAND2_X1
xU9874 n6516 n7130 n7126 VDD GND NOR2_X1
xU9875 n8333 n845 n7130 VDD GND NAND2_X1
xU9876 n6418 n6698 n6694 VDD GND NOR2_X1
xU9877 n8333 n879 n6698 VDD GND NAND2_X1
xU9878 n6488 n6982 n6978 VDD GND NOR2_X1
xU9879 n8333 n857 n6982 VDD GND NAND2_X1
xU9880 n6495 n7009 n7005 VDD GND NOR2_X1
xU9881 n8333 n854 n7009 VDD GND NAND2_X1
xU9882 n6551 n7230 n7226 VDD GND NOR2_X1
xU9883 n8332 n839 n7230 VDD GND NAND2_X1
xU9884 n6607 n7456 n7447 VDD GND NOR2_X1
xU9885 n8332 n824 n7456 VDD GND NAND2_X1
xU9886 n6411 n6669 n6665 VDD GND NOR2_X1
xU9887 n8334 n880 n6669 VDD GND NAND2_X1
xU9888 n6544 n7201 n7197 VDD GND NOR2_X1
xU9889 n8333 n840 n7201 VDD GND NAND2_X1
xU9890 n5293 n832 n5292 VDD GND NOR2_X1
xU9891 n5294 n5295 n5293 VDD GND NOR2_X1
xU9892 n8432 n370 n5295 VDD GND NOR2_X1
xU9893 n8398 n5297 n5294 VDD GND NOR2_X1
xU9894 n6904 n865 n6903 VDD GND NOR2_X1
xU9895 n6905 n8296 n6904 VDD GND NOR2_X1
xU9896 n6460 n8338 n6905 VDD GND AND2_X1
xU9897 n7348 n830 n7347 VDD GND NOR2_X1
xU9898 n7349 n8304 n7348 VDD GND NOR2_X1
xU9899 n6572 n8339 n7349 VDD GND AND2_X1
xU9900 n6667 n880 n6666 VDD GND NOR2_X1
xU9901 n6668 n8292 n6667 VDD GND NOR2_X1
xU9902 n6411 n8338 n6668 VDD GND AND2_X1
xU9903 n7449 n824 n7448 VDD GND NOR2_X1
xU9904 n7450 n8306 n7449 VDD GND NOR2_X1
xU9905 n6607 n8334 n7450 VDD GND AND2_X1
xU9906 \AES_Comp_ENCa/KrgX_9 n7018 n6966 VDD GND NAND2_X1
xU9907 n5736 n5708 n5715 VDD GND NAND2_X1
xU9908 \AES_Comp_ENCa/KrgX_22 n6858 n6818 VDD GND NAND2_X1
xU9909 n3310 n3366 n3350 VDD GND NAND2_X1
xU9910 n7428 n825 n7427 VDD GND NOR2_X1
xU9911 n7429 n8306 n7428 VDD GND NOR2_X1
xU9912 n6600 n8339 n7429 VDD GND AND2_X1
xU9913 n7336 n831 n7335 VDD GND NOR2_X1
xU9914 n7337 n8303 n7336 VDD GND NOR2_X1
xU9915 n6565 n8339 n7337 VDD GND AND2_X1
xU9916 n6892 n866 n6891 VDD GND NOR2_X1
xU9917 n6893 n8295 n6892 VDD GND NOR2_X1
xU9918 n6453 n8338 n6893 VDD GND AND2_X1
xU9919 n7128 n845 n7127 VDD GND NOR2_X1
xU9920 n7129 n8300 n7128 VDD GND NOR2_X1
xU9921 n6516 n8339 n7129 VDD GND AND2_X1
xU9922 n5460 n826 n5459 VDD GND NOR2_X1
xU9923 n5461 n5462 n5460 VDD GND NOR2_X1
xU9924 n8433 n5463 n5462 VDD GND NOR2_X1
xU9925 n8398 n347 n5461 VDD GND NOR2_X1
xU9926 n7398 n826 n7397 VDD GND NOR2_X1
xU9927 n7399 n8305 n7398 VDD GND NOR2_X1
xU9928 n8329 n6593 n7399 VDD GND NOR2_X1
xU9929 n2731 n928 n2730 VDD GND NOR2_X1
xU9930 n2732 n2733 n2731 VDD GND NOR2_X1
xU9931 n8427 n203 n2733 VDD GND NOR2_X1
xU9932 n8392 n2734 n2732 VDD GND NOR2_X1
xU9933 Dout_E_73 n5689 n5564 VDD GND NAND2_X1
xU9934 n5441 n827 n5440 VDD GND NOR2_X1
xU9935 n5442 n5443 n5441 VDD GND NOR2_X1
xU9936 n8432 n5013 n5443 VDD GND NOR2_X1
xU9937 n8398 n5444 n5442 VDD GND NOR2_X1
xU9938 n3067 n3274 n3267 VDD GND NAND2_X1
xU9939 n1820 n2113 n2101 VDD GND NAND2_X1
xU9940 n5848 n5607 n5823 VDD GND NAND2_X1
xU9941 n4804 n879 n4803 VDD GND NOR2_X1
xU9942 n4805 n4806 n4804 VDD GND NOR2_X1
xU9943 n8431 n343 n4806 VDD GND NOR2_X1
xU9944 n8396 n4807 n4805 VDD GND NOR2_X1
xU9945 \AES_Comp_ENCa/KrgX_121 n1143 n1137 VDD GND NOR2_X1
xU9946 n1144 n1145 n1143 VDD GND NOR2_X1
xU9947 n8425 n1146 n1145 VDD GND NOR2_X1
xU9948 n8390 n1142 n1144 VDD GND NOR2_X1
xU9949 n2528 n936 n2527 VDD GND NOR2_X1
xU9950 n2529 n2530 n2528 VDD GND NOR2_X1
xU9951 n8426 n421 n2530 VDD GND NOR2_X1
xU9952 n8392 n2531 n2529 VDD GND NOR2_X1
xU9953 \AES_Comp_ENCa/KrgX_78 n2655 n2648 VDD GND NOR2_X1
xU9954 n2656 n2657 n2655 VDD GND NOR2_X1
xU9955 n8427 n2653 n2657 VDD GND NOR2_X1
xU9956 n8392 n2654 n2656 VDD GND NOR2_X1
xU9957 \AES_Comp_ENCa/KrgX_33 n4306 n4300 VDD GND NOR2_X1
xU9958 n4307 n4308 n4306 VDD GND NOR2_X1
xU9959 n8430 n470 n4308 VDD GND NOR2_X1
xU9960 n8396 n4305 n4307 VDD GND NOR2_X1
xU9961 n3468 n916 n3467 VDD GND NOR2_X1
xU9962 n3469 n3470 n3468 VDD GND NOR2_X1
xU9963 n8428 n448 n3470 VDD GND NOR2_X1
xU9964 n8393 n3472 n3469 VDD GND NOR2_X1
xU9965 n4903 n867 n4902 VDD GND NOR2_X1
xU9966 n4904 n4905 n4903 VDD GND NOR2_X1
xU9967 n8431 n633 n4905 VDD GND NOR2_X1
xU9968 n8396 n4907 n4904 VDD GND NOR2_X1
xU9969 \AES_Comp_ENCa/KrgX_38 n4092 n4085 VDD GND NOR2_X1
xU9970 n4093 n4094 n4092 VDD GND NOR2_X1
xU9971 n8430 n4090 n4094 VDD GND NOR2_X1
xU9972 n8395 n4091 n4093 VDD GND NOR2_X1
xU9973 n2322 n944 n2321 VDD GND NOR2_X1
xU9974 n2323 n2324 n2322 VDD GND NOR2_X1
xU9975 n8425 n548 n2324 VDD GND NOR2_X1
xU9976 n8390 n2326 n2323 VDD GND NOR2_X1
xU9977 \AES_Comp_ENCa/KrgX_118 n1213 n1207 VDD GND NOR2_X1
xU9978 n1214 n1215 n1213 VDD GND NOR2_X1
xU9979 n8424 n1201 n1215 VDD GND NOR2_X1
xU9980 n8389 n1212 n1214 VDD GND NOR2_X1
xU9981 n2434 n940 n2433 VDD GND NOR2_X1
xU9982 n2435 n2436 n2434 VDD GND NOR2_X1
xU9983 n8426 n423 n2436 VDD GND NOR2_X1
xU9984 n8391 n2438 n2435 VDD GND NOR2_X1
xU9985 n4217 n888 n4216 VDD GND NOR2_X1
xU9986 n4218 n4219 n4217 VDD GND NOR2_X1
xU9987 n8430 n3776 n4219 VDD GND NOR2_X1
xU9988 n8395 n4220 n4218 VDD GND NOR2_X1
xU9989 n2975 n920 n2974 VDD GND NOR2_X1
xU9990 n2976 n2977 n2975 VDD GND NOR2_X1
xU9991 n8428 n2978 n2977 VDD GND NOR2_X1
xU9992 n8393 n2979 n2976 VDD GND NOR2_X1
xU9993 \AES_Comp_ENCa/KrgX_85 n2484 n2477 VDD GND NOR2_X1
xU9994 n2485 n2486 n2484 VDD GND NOR2_X1
xU9995 n8426 n424 n2486 VDD GND NOR2_X1
xU9996 n8392 n2483 n2485 VDD GND NOR2_X1
xU9997 \AES_Comp_ENCa/KrgX_41 n4017 n4010 VDD GND NOR2_X1
xU9998 n4018 n4019 n4017 VDD GND NOR2_X1
xU9999 n8430 n604 n4019 VDD GND NOR2_X1
xU10000 n8395 n4016 n4018 VDD GND NOR2_X1
xU10001 n1058 n977 n1057 VDD GND NOR2_X1
xU10002 n1059 n1060 n1058 VDD GND NOR2_X1
xU10003 n8425 n1061 n1060 VDD GND NOR2_X1
xU10004 n8391 n1062 n1059 VDD GND NOR2_X1
xU10005 n5161 n844 n5160 VDD GND NOR2_X1
xU10006 n5162 n5163 n5161 VDD GND NOR2_X1
xU10007 n8432 n504 n5163 VDD GND NOR2_X1
xU10008 n8397 n5165 n5162 VDD GND NOR2_X1
xU10009 \AES_Comp_ENCa/KrgX_102 n1606 n1599 VDD GND NOR2_X1
xU10010 n1607 n1608 n1606 VDD GND NOR2_X1
xU10011 n8424 n1604 n1608 VDD GND NOR2_X1
xU10012 n8389 n1605 n1607 VDD GND NOR2_X1
xU10013 n1500 n959 n1499 VDD GND NOR2_X1
xU10014 n1501 n1502 n1500 VDD GND NOR2_X1
xU10015 n8424 n401 n1502 VDD GND NOR2_X1
xU10016 n8390 n1504 n1501 VDD GND NOR2_X1
xU10017 \AES_Comp_ENCa/KrgX_80 n2610 n2603 VDD GND NOR2_X1
xU10018 n2611 n2612 n2610 VDD GND NOR2_X1
xU10019 n8427 n419 n2612 VDD GND NOR2_X1
xU10020 n8392 n2609 n2611 VDD GND NOR2_X1
xU10021 n1111 n975 n1110 VDD GND NOR2_X1
xU10022 n1112 n1113 n1111 VDD GND NOR2_X1
xU10023 n8425 n1114 n1113 VDD GND NOR2_X1
xU10024 n8391 n1115 n1112 VDD GND NOR2_X1
xU10025 \AES_Comp_ENCa/KrgX_89 n2381 n2375 VDD GND NOR2_X1
xU10026 n2382 n2383 n2381 VDD GND NOR2_X1
xU10027 n8426 n2384 n2383 VDD GND NOR2_X1
xU10028 n8391 n2380 n2382 VDD GND NOR2_X1
xU10029 n1086 n976 n1085 VDD GND NOR2_X1
xU10030 n1087 n1088 n1086 VDD GND NOR2_X1
xU10031 n8425 n1089 n1088 VDD GND NOR2_X1
xU10032 n8390 n1090 n1087 VDD GND NOR2_X1
xU10033 n2349 n943 n2348 VDD GND NOR2_X1
xU10034 n2350 n2351 n2349 VDD GND NOR2_X1
xU10035 n8425 n553 n2351 VDD GND NOR2_X1
xU10036 n8391 n2353 n2350 VDD GND NOR2_X1
xU10037 \AES_Comp_ENCa/KrgX_70 n2853 n2847 VDD GND NOR2_X1
xU10038 n2854 n2855 n2853 VDD GND NOR2_X1
xU10039 n8427 n585 n2855 VDD GND NOR2_X1
xU10040 n8393 n2852 n2854 VDD GND NOR2_X1
xU10041 \AES_Comp_ENCa/KrgX_110 n1407 n1400 VDD GND NOR2_X1
xU10042 n1408 n1409 n1407 VDD GND NOR2_X1
xU10043 n8423 n403 n1409 VDD GND NOR2_X1
xU10044 n8388 n1406 n1408 VDD GND NOR2_X1
xU10045 n2827 n924 n2826 VDD GND NOR2_X1
xU10046 n2828 n2829 n2827 VDD GND NOR2_X1
xU10047 n8427 n575 n2829 VDD GND NOR2_X1
xU10048 n8393 n2831 n2828 VDD GND NOR2_X1
xU10049 \AES_Comp_ENCa/KrgX_25 n4863 n4856 VDD GND NOR2_X1
xU10050 n4864 n4865 n4863 VDD GND NOR2_X1
xU10051 n8431 n320 n4865 VDD GND NOR2_X1
xU10052 n8396 n4862 n4864 VDD GND NOR2_X1
xU10053 n986 n980 n985 VDD GND NOR2_X1
xU10054 n987 n988 n986 VDD GND NOR2_X1
xU10055 n8426 n990 n988 VDD GND NOR2_X1
xU10056 n8391 n992 n987 VDD GND NOR2_X1
xU10057 \AES_Comp_ENCa/KrgX_57 n3627 n3620 VDD GND NOR2_X1
xU10058 n3628 n3629 n3627 VDD GND NOR2_X1
xU10059 n8428 n446 n3629 VDD GND NOR2_X1
xU10060 n8394 n3626 n3628 VDD GND NOR2_X1
xU10061 n3667 n908 n3666 VDD GND NOR2_X1
xU10062 n3668 n3669 n3667 VDD GND NOR2_X1
xU10063 n8428 n281 n3669 VDD GND NOR2_X1
xU10064 n8394 n3671 n3668 VDD GND NOR2_X1
xU10065 \AES_Comp_ENCa/KrgX_9 n5244 n5238 VDD GND NOR2_X1
xU10066 n5245 n5246 n5244 VDD GND NOR2_X1
xU10067 n8432 n5247 n5246 VDD GND NOR2_X1
xU10068 n8397 n5243 n5245 VDD GND NOR2_X1
xU10069 n3594 n911 n3593 VDD GND NOR2_X1
xU10070 n3595 n3596 n3594 VDD GND NOR2_X1
xU10071 n8428 n444 n3596 VDD GND NOR2_X1
xU10072 n8394 n3598 n3595 VDD GND NOR2_X1
xU10073 \AES_Comp_ENCa/KrgX_48 n3849 n3842 VDD GND NOR2_X1
xU10074 n3850 n3851 n3849 VDD GND NOR2_X1
xU10075 n8429 n257 n3851 VDD GND NOR2_X1
xU10076 n8394 n3848 n3850 VDD GND NOR2_X1
xU10077 \AES_Comp_ENCa/KrgX_17 n5050 n5044 VDD GND NOR2_X1
xU10078 n5051 n5052 n5050 VDD GND NOR2_X1
xU10079 n8431 n5033 n5052 VDD GND NOR2_X1
xU10080 n8397 n5049 n5051 VDD GND NOR2_X1
xU10081 n5368 n829 n5367 VDD GND NOR2_X1
xU10082 n5369 n5370 n5368 VDD GND NOR2_X1
xU10083 n8432 n4795 n5370 VDD GND NOR2_X1
xU10084 n8398 n346 n5369 VDD GND NOR2_X1
xU10085 n7540 n7541 n7505 VDD GND NAND2_X1
xU10086 n7437 n7521 n7540 VDD GND OR2_X1
xU10087 n7437 \AES_Comp_ENCa/KrgX_25 n7541 VDD GND NAND2_X1
xU10088 n8331 n7141 n7137 VDD GND NOR2_X1
xU10089 n6523 n844 n7141 VDD GND NAND2_X1
xU10090 n8331 n7388 n7384 VDD GND NOR2_X1
xU10091 n6586 n827 n7388 VDD GND NAND2_X1
xU10092 n8330 n6940 n6936 VDD GND NOR2_X1
xU10093 n6474 n861 n6940 VDD GND NAND2_X1
xU10094 \AES_Comp_ENCa/KrgX_14 n7074 n7048 VDD GND NAND2_X1
xU10095 n2807 n925 n2806 VDD GND NOR2_X1
xU10096 n2808 n2809 n2807 VDD GND NOR2_X1
xU10097 n2426 n8411 n2809 VDD GND NOR2_X1
xU10098 n2810 n8379 n2808 VDD GND NOR2_X1
xU10099 n3911 n898 n3910 VDD GND NOR2_X1
xU10100 n3912 n3913 n3911 VDD GND NOR2_X1
xU10101 n3528 n8407 n3913 VDD GND NOR2_X1
xU10102 n3914 n8382 n3912 VDD GND NOR2_X1
xU10103 \AES_Comp_ENCa/KrgX_19 n5003 n4997 VDD GND NOR2_X1
xU10104 n5004 n5005 n5003 VDD GND NOR2_X1
xU10105 n630 n8404 n5005 VDD GND NOR2_X1
xU10106 n5002 n8386 n5004 VDD GND NOR2_X1
xU10107 \AES_Comp_ENCa/KrgX_18 n5027 n5020 VDD GND NOR2_X1
xU10108 n5028 n5029 n5027 VDD GND NOR2_X1
xU10109 n5025 n8404 n5029 VDD GND NOR2_X1
xU10110 n5026 n8386 n5028 VDD GND NOR2_X1
xU10111 \AES_Comp_ENCa/KrgX_52 n3741 n3734 VDD GND NOR2_X1
xU10112 n3742 n3743 n3741 VDD GND NOR2_X1
xU10113 n290 n8408 n3743 VDD GND NOR2_X1
xU10114 n3740 n8382 n3742 VDD GND NOR2_X1
xU10115 \AES_Comp_ENCa/KrgX_44 n3935 n3929 VDD GND NOR2_X1
xU10116 n3936 n3937 n3935 VDD GND NOR2_X1
xU10117 n607 n8407 n3937 VDD GND NOR2_X1
xU10118 n3934 n8383 n3936 VDD GND NOR2_X1
xU10119 \AES_Comp_ENCa/KrgX_79 n2631 n2625 VDD GND NOR2_X1
xU10120 n2632 n2633 n2631 VDD GND NOR2_X1
xU10121 n2634 n8412 n2633 VDD GND NOR2_X1
xU10122 n2630 n8378 n2632 VDD GND NOR2_X1
xU10123 n3690 n907 n3689 VDD GND NOR2_X1
xU10124 n3691 n3692 n3690 VDD GND NOR2_X1
xU10125 n3693 n8408 n3692 VDD GND NOR2_X1
xU10126 n3694 n8381 n3691 VDD GND NOR2_X1
xU10127 n4950 n865 n4949 VDD GND NOR2_X1
xU10128 n4951 n4952 n4950 VDD GND NOR2_X1
xU10129 n631 n8404 n4952 VDD GND NOR2_X1
xU10130 n4953 n8385 n4951 VDD GND NOR2_X1
xU10131 \AES_Comp_ENCa/KrgX_103 n1584 n1577 VDD GND NOR2_X1
xU10132 n1585 n1586 n1584 VDD GND NOR2_X1
xU10133 n1582 n8408 n1586 VDD GND NOR2_X1
xU10134 n1583 n8382 n1585 VDD GND NOR2_X1
xU10135 n1233 n970 n1232 VDD GND NOR2_X1
xU10136 n1234 n1235 n1233 VDD GND NOR2_X1
xU10137 n523 n8404 n1235 VDD GND NOR2_X1
xU10138 n1236 n8385 n1234 VDD GND NOR2_X1
xU10139 n4758 n882 n4757 VDD GND NOR2_X1
xU10140 n4759 n4760 n4758 VDD GND NOR2_X1
xU10141 n4745 n8405 n4760 VDD GND NOR2_X1
xU10142 n4761 n8385 n4759 VDD GND NOR2_X1
xU10143 \AES_Comp_ENCa/KrgX_36 n4149 n4142 VDD GND NOR2_X1
xU10144 n4150 n4151 n4149 VDD GND NOR2_X1
xU10145 n4147 n8406 n4151 VDD GND NOR2_X1
xU10146 n4148 n8384 n4150 VDD GND NOR2_X1
xU10147 \AES_Comp_ENCa/KrgX_11 n5197 n5191 VDD GND NOR2_X1
xU10148 n5198 n5199 n5197 VDD GND NOR2_X1
xU10149 n497 n8403 n5199 VDD GND NOR2_X1
xU10150 n5196 n8386 n5198 VDD GND NOR2_X1
xU10151 \AES_Comp_ENCa/KrgX_107 n1482 n1475 VDD GND NOR2_X1
xU10152 n1483 n1484 n1482 VDD GND NOR2_X1
xU10153 n397 n8407 n1484 VDD GND NOR2_X1
xU10154 n1481 n8383 n1483 VDD GND NOR2_X1
xU10155 n1037 n978 n1036 VDD GND NOR2_X1
xU10156 n1038 n1039 n1037 VDD GND NOR2_X1
xU10157 n1040 n8402 n1039 VDD GND NOR2_X1
xU10158 n1041 n8387 n1038 VDD GND NOR2_X1
xU10159 n3519 n914 n3518 VDD GND NOR2_X1
xU10160 n3520 n3521 n3519 VDD GND NOR2_X1
xU10161 n3504 n8409 n3521 VDD GND NOR2_X1
xU10162 n3522 n8380 n3520 VDD GND NOR2_X1
xU10163 n1626 n954 n1625 VDD GND NOR2_X1
xU10164 n1627 n1628 n1626 VDD GND NOR2_X1
xU10165 n161 n8408 n1628 VDD GND NOR2_X1
xU10166 n1629 n8381 n1627 VDD GND NOR2_X1
xU10167 n3715 n906 n3714 VDD GND NOR2_X1
xU10168 n3716 n3717 n3715 VDD GND NOR2_X1
xU10169 n269 n8408 n3717 VDD GND NOR2_X1
xU10170 n3718 n8381 n3716 VDD GND NOR2_X1
xU10171 \AES_Comp_ENCa/KrgX_28 n4783 n4777 VDD GND NOR2_X1
xU10172 n4784 n4785 n4783 VDD GND NOR2_X1
xU10173 n4771 n8405 n4785 VDD GND NOR2_X1
xU10174 n4782 n8385 n4784 VDD GND NOR2_X1
xU10175 \AES_Comp_ENCa/KrgX_92 n2299 n2292 VDD GND NOR2_X1
xU10176 n2300 n2301 n2299 VDD GND NOR2_X1
xU10177 n2297 n8411 n2301 VDD GND NOR2_X1
xU10178 n2298 n8379 n2300 VDD GND NOR2_X1
xU10179 \AES_Comp_ENCa/KrgX_108 n1451 n1445 VDD GND NOR2_X1
xU10180 n1452 n1453 n1451 VDD GND NOR2_X1
xU10181 n1072 n8406 n1453 VDD GND NOR2_X1
xU10182 n1450 n8383 n1452 VDD GND NOR2_X1
xU10183 \AES_Comp_ENCa/KrgX_51 n3765 n3758 VDD GND NOR2_X1
xU10184 n3766 n3767 n3765 VDD GND NOR2_X1
xU10185 n262 n8408 n3767 VDD GND NOR2_X1
xU10186 n3764 n8382 n3766 VDD GND NOR2_X1
xU10187 n1425 n962 n1424 VDD GND NOR2_X1
xU10188 n1426 n1427 n1425 VDD GND NOR2_X1
xU10189 n1428 n8406 n1427 VDD GND NOR2_X1
xU10190 n1429 n8383 n1426 VDD GND NOR2_X1
xU10191 n5141 n845 n5140 VDD GND NOR2_X1
xU10192 n5142 n5143 n5141 VDD GND NOR2_X1
xU10193 n499 n8403 n5143 VDD GND NOR2_X1
xU10194 n5144 n8386 n5142 VDD GND NOR2_X1
xU10195 n1529 n958 n1528 VDD GND NOR2_X1
xU10196 n1530 n1531 n1529 VDD GND NOR2_X1
xU10197 n1515 n8407 n1531 VDD GND NOR2_X1
xU10198 n1532 n8382 n1530 VDD GND NOR2_X1
xU10199 n5042 n5043 n7956 VDD GND NAND2_X1
xU10200 n5065 n5066 n5042 VDD GND NOR2_X1
xU10201 n5044 n5045 n5043 VDD GND NOR2_X1
xU10202 n8369 n303 n5066 VDD GND NOR2_X1
xU10203 \AES_Comp_ENCa/KrgX_59 n3572 n3565 VDD GND NOR2_X1
xU10204 n3573 n3574 n3572 VDD GND NOR2_X1
xU10205 n450 n8409 n3574 VDD GND NOR2_X1
xU10206 n3571 n8381 n3573 VDD GND NOR2_X1
xU10207 \AES_Comp_ENCa/KrgX_26 n4835 n4828 VDD GND NOR2_X1
xU10208 n4836 n4837 n4835 VDD GND NOR2_X1
xU10209 n332 n8405 n4837 VDD GND NOR2_X1
xU10210 n4834 n8385 n4836 VDD GND NOR2_X1
xU10211 \AES_Comp_ENCa/KrgX_114 n1312 n1305 VDD GND NOR2_X1
xU10212 n1313 n1314 n1312 VDD GND NOR2_X1
xU10213 n527 n8405 n1314 VDD GND NOR2_X1
xU10214 n1311 n8385 n1313 VDD GND NOR2_X1
xU10215 \AES_Comp_ENCa/KrgX_99 n1731 n1725 VDD GND NOR2_X1
xU10216 n1732 n1733 n1731 VDD GND NOR2_X1
xU10217 n1734 n8409 n1733 VDD GND NOR2_X1
xU10218 n1730 n8381 n1732 VDD GND NOR2_X1
xU10219 \AES_Comp_ENCa/KrgX_76 n2704 n2698 VDD GND NOR2_X1
xU10220 n2705 n2706 n2704 VDD GND NOR2_X1
xU10221 n2311 n8411 n2706 VDD GND NOR2_X1
xU10222 n2703 n8379 n2705 VDD GND NOR2_X1
xU10223 \AES_Comp_ENCa/KrgX_2 n5465 n5458 VDD GND NOR2_X1
xU10224 n5466 n5467 n5465 VDD GND NOR2_X1
xU10225 n373 n8402 n5467 VDD GND NOR2_X1
xU10226 n5464 n8388 n5466 VDD GND NOR2_X1
xU10227 \AES_Comp_ENCa/KrgX_115 n1285 n1278 VDD GND NOR2_X1
xU10228 n1286 n1287 n1285 VDD GND NOR2_X1
xU10229 n522 n8405 n1287 VDD GND NOR2_X1
xU10230 n1284 n8385 n1286 VDD GND NOR2_X1
xU10231 \AES_Comp_ENCa/KrgX_43 n3965 n3959 VDD GND NOR2_X1
xU10232 n3966 n3967 n3965 VDD GND NOR2_X1
xU10233 n602 n8407 n3967 VDD GND NOR2_X1
xU10234 n3964 n8383 n3966 VDD GND NOR2_X1
xU10235 n3645 n909 n3644 VDD GND NOR2_X1
xU10236 n3646 n3647 n3645 VDD GND NOR2_X1
xU10237 n3648 n8409 n3647 VDD GND NOR2_X1
xU10238 n3649 n8381 n3646 VDD GND NOR2_X1
xU10239 \AES_Comp_ENCa/KrgX_84 n2507 n2501 VDD GND NOR2_X1
xU10240 n2508 n2509 n2507 VDD GND NOR2_X1
xU10241 n2510 n8412 n2509 VDD GND NOR2_X1
xU10242 n2506 n8378 n2508 VDD GND NOR2_X1
xU10243 \AES_Comp_ENCa/KrgX_116 n1259 n1252 VDD GND NOR2_X1
xU10244 n1260 n1261 n1259 VDD GND NOR2_X1
xU10245 n528 n8404 n1261 VDD GND NOR2_X1
xU10246 n1258 n8385 n1260 VDD GND NOR2_X1
xU10247 \AES_Comp_ENCa/KrgX_82 n2556 n2549 VDD GND NOR2_X1
xU10248 n2557 n2558 n2556 VDD GND NOR2_X1
xU10249 n422 n8412 n2558 VDD GND NOR2_X1
xU10250 n2555 n8378 n2557 VDD GND NOR2_X1
xU10251 n2674 n930 n2673 VDD GND NOR2_X1
xU10252 n2675 n2676 n2674 VDD GND NOR2_X1
xU10253 n217 n8411 n2676 VDD GND NOR2_X1
xU10254 n2678 n8378 n2675 VDD GND NOR2_X1
xU10255 n5583 n824 n5582 VDD GND NOR2_X1
xU10256 n5584 n5585 n5583 VDD GND NOR2_X1
xU10257 n4895 n8407 n5585 VDD GND NOR2_X1
xU10258 n5586 n8388 n5584 VDD GND NOR2_X1
xU10259 n1867 n949 n1866 VDD GND NOR2_X1
xU10260 n1868 n1869 n1867 VDD GND NOR2_X1
xU10261 n1870 n8409 n1869 VDD GND NOR2_X1
xU10262 n1871 n8380 n1868 VDD GND NOR2_X1
xU10263 n2458 n939 n2457 VDD GND NOR2_X1
xU10264 n2459 n2460 n2458 VDD GND NOR2_X1
xU10265 n2461 n8412 n2460 VDD GND NOR2_X1
xU10266 n2462 n8378 n2459 VDD GND NOR2_X1
xU10267 n4927 n866 n4926 VDD GND NOR2_X1
xU10268 n4928 n4929 n4927 VDD GND NOR2_X1
xU10269 n638 n8404 n4929 VDD GND NOR2_X1
xU10270 n4931 n8386 n4928 VDD GND NOR2_X1
xU10271 n2874 n922 n2873 VDD GND NOR2_X1
xU10272 n2875 n2876 n2874 VDD GND NOR2_X1
xU10273 n2877 n8410 n2876 VDD GND NOR2_X1
xU10274 n2878 n8379 n2875 VDD GND NOR2_X1
xU10275 n1014 n979 n1013 VDD GND NOR2_X1
xU10276 n1015 n1016 n1014 VDD GND NOR2_X1
xU10277 n663 n8402 n1016 VDD GND NOR2_X1
xU10278 n1017 n8388 n1015 VDD GND NOR2_X1
xU10279 \AES_Comp_ENCa/KrgX_20 n4978 n4971 VDD GND NOR2_X1
xU10280 n4979 n4980 n4978 VDD GND NOR2_X1
xU10281 n636 n8404 n4980 VDD GND NOR2_X1
xU10282 n4977 n8386 n4979 VDD GND NOR2_X1
xU10283 n4733 n883 n4732 VDD GND NOR2_X1
xU10284 n4734 n4735 n4733 VDD GND NOR2_X1
xU10285 n4736 n8405 n4735 VDD GND NOR2_X1
xU10286 n4737 n8384 n4734 VDD GND NOR2_X1
xU10287 \AES_Comp_ENCa/KrgX_39 n4068 n4062 VDD GND NOR2_X1
xU10288 n4069 n4070 n4068 VDD GND NOR2_X1
xU10289 n469 n8406 n4070 VDD GND NOR2_X1
xU10290 n4067 n8383 n4069 VDD GND NOR2_X1
xU10291 \AES_Comp_ENCa/KrgX_60 n3545 n3539 VDD GND NOR2_X1
xU10292 n3546 n3547 n3545 VDD GND NOR2_X1
xU10293 n449 n8409 n3547 VDD GND NOR2_X1
xU10294 n3544 n8381 n3546 VDD GND NOR2_X1
xU10295 \AES_Comp_ENCa/KrgX_10 n5220 n5213 VDD GND NOR2_X1
xU10296 n5221 n5222 n5220 VDD GND NOR2_X1
xU10297 n5218 n8403 n5222 VDD GND NOR2_X1
xU10298 n5219 n8387 n5221 VDD GND NOR2_X1
xU10299 \AES_Comp_ENCa/KrgX_111 n1383 n1376 VDD GND NOR2_X1
xU10300 n1384 n1385 n1383 VDD GND NOR2_X1
xU10301 n1381 n8406 n1385 VDD GND NOR2_X1
xU10302 n1382 n8384 n1384 VDD GND NOR2_X1
xU10303 n5315 n831 n5314 VDD GND NOR2_X1
xU10304 n5316 n5317 n5315 VDD GND NOR2_X1
xU10305 n5318 n8402 n5317 VDD GND NOR2_X1
xU10306 n5319 n8388 n5316 VDD GND NOR2_X1
xU10307 \AES_Comp_ENCa/KrgX_50 n3790 n3783 VDD GND NOR2_X1
xU10308 n3791 n3792 n3790 VDD GND NOR2_X1
xU10309 n284 n8408 n3792 VDD GND NOR2_X1
xU10310 n3789 n8382 n3791 VDD GND NOR2_X1
xU10311 n3494 n915 n3493 VDD GND NOR2_X1
xU10312 n3495 n3496 n3494 VDD GND NOR2_X1
xU10313 n453 n8409 n3496 VDD GND NOR2_X1
xU10314 n3497 n8380 n3495 VDD GND NOR2_X1
xU10315 n2408 n941 n2407 VDD GND NOR2_X1
xU10316 n2409 n2410 n2408 VDD GND NOR2_X1
xU10317 n2411 n8411 n2410 VDD GND NOR2_X1
xU10318 n2412 n8378 n2409 VDD GND NOR2_X1
xU10319 \AES_Comp_ENCa/KrgX_100 n1660 n1654 VDD GND NOR2_X1
xU10320 n1661 n1662 n1660 VDD GND NOR2_X1
xU10321 n166 n8409 n1662 VDD GND NOR2_X1
xU10322 n1659 n8381 n1661 VDD GND NOR2_X1
xU10323 \AES_Comp_ENCa/KrgX_31 n4708 n4701 VDD GND NOR2_X1
xU10324 n4709 n4710 n4708 VDD GND NOR2_X1
xU10325 n328 n8405 n4710 VDD GND NOR2_X1
xU10326 n4707 n8384 n4709 VDD GND NOR2_X1
xU10327 \AES_Comp_ENCa/KrgX_42 n3991 n3984 VDD GND NOR2_X1
xU10328 n3992 n3993 n3991 VDD GND NOR2_X1
xU10329 n3989 n8407 n3993 VDD GND NOR2_X1
xU10330 n3990 n8384 n3992 VDD GND NOR2_X1
xU10331 \AES_Comp_ENCa/KrgX_68 n2907 n2901 VDD GND NOR2_X1
xU10332 n2908 n2909 n2907 VDD GND NOR2_X1
xU10333 n2313 n8410 n2909 VDD GND NOR2_X1
xU10334 n2906 n8380 n2908 VDD GND NOR2_X1
xU10335 n5117 n846 n5116 VDD GND NOR2_X1
xU10336 n5118 n5119 n5117 VDD GND NOR2_X1
xU10337 n5120 n8403 n5119 VDD GND NOR2_X1
xU10338 n5121 n8387 n5118 VDD GND NOR2_X1
xU10339 n5072 n854 n5071 VDD GND NOR2_X1
xU10340 n5073 n5074 n5072 VDD GND NOR2_X1
xU10341 n5075 n8404 n5074 VDD GND NOR2_X1
xU10342 n5076 n8386 n5073 VDD GND NOR2_X1
xU10343 n5266 n5267 n7965 VDD GND NAND2_X1
xU10344 n5286 n5287 n5266 VDD GND NOR2_X1
xU10345 n5268 n5269 n5267 VDD GND NOR2_X1
xU10346 n8370 n243 n5287 VDD GND NOR2_X1
xU10347 n4347 n885 n4346 VDD GND NOR2_X1
xU10348 n4348 n4349 n4347 VDD GND NOR2_X1
xU10349 n3856 n8406 n4349 VDD GND NOR2_X1
xU10350 n4350 n8384 n4348 VDD GND NOR2_X1
xU10351 \AES_Comp_ENCa/KrgX_66 n3001 n2994 VDD GND NOR2_X1
xU10352 n3002 n3003 n3001 VDD GND NOR2_X1
xU10353 n2999 n8412 n3003 VDD GND NOR2_X1
xU10354 n3000 n8380 n3002 VDD GND NOR2_X1
xU10355 \AES_Comp_ENCa/KrgX_74 n2761 n2754 VDD GND NOR2_X1
xU10356 n2762 n2763 n2761 VDD GND NOR2_X1
xU10357 n206 n8411 n2763 VDD GND NOR2_X1
xU10358 n2760 n8379 n2762 VDD GND NOR2_X1
xU10359 n1163 n973 n1162 VDD GND NOR2_X1
xU10360 n1164 n1165 n1163 VDD GND NOR2_X1
xU10361 n1166 n8403 n1165 VDD GND NOR2_X1
xU10362 n1167 n8387 n1164 VDD GND NOR2_X1
xU10363 \AES_Comp_ENCa/KrgX_98 n1753 n1746 VDD GND NOR2_X1
xU10364 n1754 n1755 n1753 VDD GND NOR2_X1
xU10365 n141 n8409 n1755 VDD GND NOR2_X1
xU10366 n1752 n8381 n1754 VDD GND NOR2_X1
xU10367 n4899 n4900 n7950 VDD GND NAND2_X1
xU10368 n4920 n4921 n4899 VDD GND NOR2_X1
xU10369 n4901 n4902 n4900 VDD GND NOR2_X1
xU10370 n8368 n312 n4921 VDD GND NOR2_X1
xU10371 n4969 n4970 n7953 VDD GND NAND2_X1
xU10372 n4992 n4993 n4969 VDD GND NOR2_X1
xU10373 n4971 n4972 n4970 VDD GND NOR2_X1
xU10374 n8369 n309 n4993 VDD GND NOR2_X1
xU10375 n4699 n4700 n7942 VDD GND NAND2_X1
xU10376 n4726 n4727 n4699 VDD GND NOR2_X1
xU10377 n4701 n4702 n4700 VDD GND NOR2_X1
xU10378 n8368 n369 n4727 VDD GND NOR2_X1
xU10379 n2780 n926 n2779 VDD GND NOR2_X1
xU10380 n2781 n2782 n2780 VDD GND NOR2_X1
xU10381 n234 n8411 n2782 VDD GND NOR2_X1
xU10382 n2784 n8379 n2781 VDD GND NOR2_X1
xU10383 n4826 n4827 n7947 VDD GND NAND2_X1
xU10384 n4851 n4852 n4826 VDD GND NOR2_X1
xU10385 n4828 n4829 n4827 VDD GND NOR2_X1
xU10386 n8368 n364 n4852 VDD GND NOR2_X1
xU10387 n4879 n4880 n7949 VDD GND NAND2_X1
xU10388 n4896 n4897 n4879 VDD GND NOR2_X1
xU10389 n4881 n4882 n4880 VDD GND NOR2_X1
xU10390 n8368 n361 n4897 VDD GND NOR2_X1
xU10391 n5018 n5019 n7955 VDD GND NAND2_X1
xU10392 n5039 n5040 n5018 VDD GND NOR2_X1
xU10393 n5020 n5021 n5019 VDD GND NOR2_X1
xU10394 n8369 n306 n5040 VDD GND NOR2_X1
xU10395 n5068 n5069 n7957 VDD GND NAND2_X1
xU10396 n5087 n5088 n5068 VDD GND NOR2_X1
xU10397 n5070 n5071 n5069 VDD GND NOR2_X1
xU10398 n8369 n301 n5088 VDD GND NOR2_X1
xU10399 \AES_Comp_ENCa/KrgX_47 n3869 n3862 VDD GND NOR2_X1
xU10400 n3870 n3871 n3869 VDD GND NOR2_X1
xU10401 n605 n8408 n3871 VDD GND NOR2_X1
xU10402 n3868 n8382 n3870 VDD GND NOR2_X1
xU10403 n2245 n947 n2244 VDD GND NOR2_X1
xU10404 n2246 n2247 n2245 VDD GND NOR2_X1
xU10405 n2248 n8410 n2247 VDD GND NOR2_X1
xU10406 n2249 n8380 n2246 VDD GND NOR2_X1
xU10407 n5236 n5237 n7964 VDD GND NAND2_X1
xU10408 n5263 n5264 n5236 VDD GND NOR2_X1
xU10409 n5238 n5239 n5237 VDD GND NOR2_X1
xU10410 n8370 n245 n5264 VDD GND NOR2_X1
xU10411 \AES_Comp_ENCa/KrgX_15 n5099 n5092 VDD GND NOR2_X1
xU10412 n5100 n5101 n5099 VDD GND NOR2_X1
xU10413 n501 n8403 n5101 VDD GND NOR2_X1
xU10414 n5098 n8387 n5100 VDD GND NOR2_X1
xU10415 n3058 n918 n3057 VDD GND NOR2_X1
xU10416 n3059 n3060 n3058 VDD GND NOR2_X1
xU10417 n3061 n8410 n3060 VDD GND NOR2_X1
xU10418 n3062 n8380 n3059 VDD GND NOR2_X1
xU10419 n1557 n957 n1556 VDD GND NOR2_X1
xU10420 n1558 n1559 n1557 VDD GND NOR2_X1
xU10421 n1560 n8407 n1559 VDD GND NOR2_X1
xU10422 n1561 n8382 n1558 VDD GND NOR2_X1
xU10423 n2270 n946 n2269 VDD GND NOR2_X1
xU10424 n2271 n2272 n2270 VDD GND NOR2_X1
xU10425 n549 n8410 n2272 VDD GND NOR2_X1
xU10426 n2273 n8379 n2271 VDD GND NOR2_X1
xU10427 n5339 n830 n5338 VDD GND NOR2_X1
xU10428 n5340 n5341 n5339 VDD GND NOR2_X1
xU10429 n4960 n8402 n5341 VDD GND NOR2_X1
xU10430 n5342 n8388 n5340 VDD GND NOR2_X1
xU10431 n5270 n839 n5269 VDD GND NOR2_X1
xU10432 n5271 n5272 n5270 VDD GND NOR2_X1
xU10433 n5273 n8403 n5272 VDD GND NOR2_X1
xU10434 n5274 n8387 n5271 VDD GND NOR2_X1
xU10435 n4114 n890 n4113 VDD GND NOR2_X1
xU10436 n4115 n4116 n4114 VDD GND NOR2_X1
xU10437 n471 n8406 n4116 VDD GND NOR2_X1
xU10438 n4117 n8383 n4115 VDD GND NOR2_X1
xU10439 \AES_Comp_ENCa/KrgX_119 n1188 n1181 VDD GND NOR2_X1
xU10440 n1189 n1190 n1188 VDD GND NOR2_X1
xU10441 n1186 n8404 n1190 VDD GND NOR2_X1
xU10442 n1187 n8386 n1189 VDD GND NOR2_X1
xU10443 n4043 n893 n4042 VDD GND NOR2_X1
xU10444 n4044 n4045 n4043 VDD GND NOR2_X1
xU10445 n4046 n8407 n4045 VDD GND NOR2_X1
xU10446 n4047 n8383 n4044 VDD GND NOR2_X1
xU10447 n1359 n965 n1358 VDD GND NOR2_X1
xU10448 n1360 n1361 n1359 VDD GND NOR2_X1
xU10449 n1362 n8405 n1361 VDD GND NOR2_X1
xU10450 n1363 n8384 n1360 VDD GND NOR2_X1
xU10451 \AES_Comp_ENCa/KrgX_95 n2226 n2219 VDD GND NOR2_X1
xU10452 n2227 n2228 n2226 VDD GND NOR2_X1
xU10453 n2224 n8410 n2228 VDD GND NOR2_X1
xU10454 n2225 n8380 n2227 VDD GND NOR2_X1
xU10455 n3888 n899 n3887 VDD GND NOR2_X1
xU10456 n3889 n3890 n3888 VDD GND NOR2_X1
xU10457 n610 n8407 n3890 VDD GND NOR2_X1
xU10458 n3891 n8382 n3889 VDD GND NOR2_X1
xU10459 n1332 n966 n1331 VDD GND NOR2_X1
xU10460 n1333 n1334 n1332 VDD GND NOR2_X1
xU10461 n1335 n8405 n1334 VDD GND NOR2_X1
xU10462 n1336 n8384 n1333 VDD GND NOR2_X1
xU10463 \AES_Comp_ENCa/KrgX_4 n5372 n5366 VDD GND NOR2_X1
xU10464 n5373 n5374 n5372 VDD GND NOR2_X1
xU10465 n377 n8402 n5374 VDD GND NOR2_X1
xU10466 n5371 n8388 n5373 VDD GND NOR2_X1
xU10467 n4883 n875 n4882 VDD GND NOR2_X1
xU10468 n4884 n4885 n4883 VDD GND NOR2_X1
xU10469 n4886 n8405 n4885 VDD GND NOR2_X1
xU10470 n4887 n8385 n4884 VDD GND NOR2_X1
xU10471 n3816 n902 n3815 VDD GND NOR2_X1
xU10472 n3817 n3818 n3816 VDD GND NOR2_X1
xU10473 n3819 n8408 n3818 VDD GND NOR2_X1
xU10474 n3820 n8382 n3817 VDD GND NOR2_X1
xU10475 n2577 n934 n2576 VDD GND NOR2_X1
xU10476 n2578 n2579 n2577 VDD GND NOR2_X1
xU10477 n2580 n8412 n2579 VDD GND NOR2_X1
xU10478 n2581 n8378 n2578 VDD GND NOR2_X1
xU10479 n3113 n917 n3112 VDD GND NOR2_X1
xU10480 n3114 n3115 n3113 VDD GND NOR2_X1
xU10481 n578 n8410 n3115 VDD GND NOR2_X1
xU10482 n3116 n8380 n3114 VDD GND NOR2_X1
xU10483 n1812 n950 n1811 VDD GND NOR2_X1
xU10484 n1813 n1814 n1812 VDD GND NOR2_X1
xU10485 n1815 n8409 n1814 VDD GND NOR2_X1
xU10486 n1816 n8380 n1813 VDD GND NOR2_X1
xU10487 n4729 n4730 n7943 VDD GND NAND2_X1
xU10488 n4751 n4752 n4729 VDD GND NOR2_X1
xU10489 n4731 n4732 n4730 VDD GND NOR2_X1
xU10490 n8368 n368 n4752 VDD GND NOR2_X1
xU10491 n5335 n5336 n7968 VDD GND NAND2_X1
xU10492 n5361 n5362 n5335 VDD GND NOR2_X1
xU10493 n5337 n5338 n5336 VDD GND NOR2_X1
xU10494 n195 n8357 n5362 VDD GND NOR2_X1
xU10495 n5090 n5091 n7958 VDD GND NAND2_X1
xU10496 n5110 n5111 n5090 VDD GND NOR2_X1
xU10497 n5092 n5093 n5091 VDD GND NOR2_X1
xU10498 n8369 n255 n5111 VDD GND NOR2_X1
xU10499 n4946 n4947 n7952 VDD GND NAND2_X1
xU10500 n4966 n4967 n4946 VDD GND NOR2_X1
xU10501 n4948 n4949 n4947 VDD GND NOR2_X1
xU10502 n8369 n310 n4967 VDD GND NOR2_X1
xU10503 n4775 n4776 n7945 VDD GND NAND2_X1
xU10504 n4797 n4798 n4775 VDD GND NOR2_X1
xU10505 n4777 n4778 n4776 VDD GND NOR2_X1
xU10506 n8368 n366 n4798 VDD GND NOR2_X1
xU10507 n5289 n5290 n7966 VDD GND NAND2_X1
xU10508 n5308 n5309 n5289 VDD GND NOR2_X1
xU10509 n5291 n5292 n5290 VDD GND NOR2_X1
xU10510 n197 n8358 n5309 VDD GND NOR2_X1
xU10511 n5211 n5212 n7963 VDD GND NAND2_X1
xU10512 n5233 n5234 n5211 VDD GND NOR2_X1
xU10513 n5213 n5214 n5212 VDD GND NOR2_X1
xU10514 n8370 n248 n5234 VDD GND NOR2_X1
xU10515 n5364 n5365 n7969 VDD GND NAND2_X1
xU10516 n5434 n5435 n5364 VDD GND NOR2_X1
xU10517 n5366 n5367 n5365 VDD GND NOR2_X1
xU10518 n194 n8357 n5435 VDD GND NOR2_X1
xU10519 n5579 n5580 n7973 VDD GND NAND2_X1
xU10520 n5932 n5933 n5579 VDD GND NOR2_X1
xU10521 n5581 n5582 n5580 VDD GND NOR2_X1
xU10522 n188 n8357 n5933 VDD GND NOR2_X1
xU10523 n4923 n4924 n7951 VDD GND NAND2_X1
xU10524 n4943 n4944 n4923 VDD GND NOR2_X1
xU10525 n4925 n4926 n4924 VDD GND NOR2_X1
xU10526 n8368 n311 n4944 VDD GND NOR2_X1
xU10527 n4754 n4755 n7944 VDD GND NAND2_X1
xU10528 n4772 n4773 n4754 VDD GND NOR2_X1
xU10529 n4756 n4757 n4755 VDD GND NOR2_X1
xU10530 n8368 n367 n4773 VDD GND NOR2_X1
xU10531 n5311 n5312 n7967 VDD GND NAND2_X1
xU10532 n5332 n5333 n5311 VDD GND NOR2_X1
xU10533 n5313 n5314 n5312 VDD GND NOR2_X1
xU10534 n196 n8357 n5333 VDD GND NOR2_X1
xU10535 n5137 n5138 n7960 VDD GND NAND2_X1
xU10536 n5154 n5155 n5137 VDD GND NOR2_X1
xU10537 n5139 n5140 n5138 VDD GND NOR2_X1
xU10538 n8369 n253 n5155 VDD GND NOR2_X1
xU10539 n5113 n5114 n7959 VDD GND NAND2_X1
xU10540 n5134 n5135 n5113 VDD GND NOR2_X1
xU10541 n5115 n5116 n5114 VDD GND NOR2_X1
xU10542 n8369 n254 n5135 VDD GND NOR2_X1
xU10543 n4800 n4801 n7946 VDD GND NAND2_X1
xU10544 n4823 n4824 n4800 VDD GND NOR2_X1
xU10545 n4802 n4803 n4801 VDD GND NOR2_X1
xU10546 n8368 n365 n4824 VDD GND NOR2_X1
xU10547 n5189 n5190 n7962 VDD GND NAND2_X1
xU10548 n5208 n5209 n5189 VDD GND NOR2_X1
xU10549 n5191 n5192 n5190 VDD GND NOR2_X1
xU10550 n8370 n249 n5209 VDD GND NOR2_X1
xU10551 n4995 n4996 n7954 VDD GND NAND2_X1
xU10552 n5015 n5016 n4995 VDD GND NOR2_X1
xU10553 n4997 n4998 n4996 VDD GND NOR2_X1
xU10554 n8369 n307 n5016 VDD GND NOR2_X1
xU10555 n5437 n5438 n7970 VDD GND NAND2_X1
xU10556 n5453 n5454 n5437 VDD GND NOR2_X1
xU10557 n5439 n5440 n5438 VDD GND NOR2_X1
xU10558 n192 n8357 n5454 VDD GND NOR2_X1
xU10559 n1622 n1623 n7872 VDD GND NAND2_X1
xU10560 n1649 n1650 n1622 VDD GND NOR2_X1
xU10561 n1624 n1625 n1623 VDD GND NOR2_X1
xU10562 n8361 n598 n1650 VDD GND NOR2_X1
xU10563 n1082 n1083 n7850 VDD GND NAND2_X1
xU10564 n1104 n1105 n1082 VDD GND NOR2_X1
xU10565 n1084 n1085 n1083 VDD GND NOR2_X1
xU10566 n674 n8358 n1105 VDD GND NOR2_X1
xU10567 n1010 n1011 n7847 VDD GND NAND2_X1
xU10568 n1030 n1031 n1010 VDD GND NOR2_X1
xU10569 n1012 n1013 n1011 VDD GND NOR2_X1
xU10570 n679 n8358 n1031 VDD GND NOR2_X1
xU10571 n1107 n1108 n7851 VDD GND NAND2_X1
xU10572 n1132 n1133 n1107 VDD GND NOR2_X1
xU10573 n1109 n1110 n1108 VDD GND NOR2_X1
xU10574 n673 n8358 n1133 VDD GND NOR2_X1
xU10575 n1553 n1554 n7869 VDD GND NAND2_X1
xU10576 n1572 n1573 n1553 VDD GND NOR2_X1
xU10577 n1555 n1556 n1554 VDD GND NOR2_X1
xU10578 n8362 n617 n1573 VDD GND NOR2_X1
xU10579 n1863 n1864 n7877 VDD GND NAND2_X1
xU10580 n2214 n2215 n1863 VDD GND NOR2_X1
xU10581 n1865 n1866 n1864 VDD GND NOR2_X1
xU10582 n8362 n591 n2215 VDD GND NOR2_X1
xU10583 n1355 n1356 n7861 VDD GND NAND2_X1
xU10584 n1371 n1372 n1355 VDD GND NOR2_X1
xU10585 n1357 n1358 n1356 VDD GND NOR2_X1
xU10586 n8363 n643 n1372 VDD GND NOR2_X1
xU10587 n1229 n1230 n7856 VDD GND NAND2_X1
xU10588 n1247 n1248 n1229 VDD GND NOR2_X1
xU10589 n1231 n1232 n1230 VDD GND NOR2_X1
xU10590 n8360 n654 n1248 VDD GND NOR2_X1
xU10591 n1808 n1809 n7876 VDD GND NAND2_X1
xU10592 n1860 n1861 n1808 VDD GND NOR2_X1
xU10593 n1810 n1811 n1809 VDD GND NOR2_X1
xU10594 n8362 n593 n1861 VDD GND NOR2_X1
xU10595 n2217 n2218 n7878 VDD GND NAND2_X1
xU10596 n2238 n2239 n2217 VDD GND NOR2_X1
xU10597 n2219 n2220 n2218 VDD GND NOR2_X1
xU10598 n8364 n572 n2239 VDD GND NOR2_X1
xU10599 n2623 n2624 n7894 VDD GND NAND2_X1
xU10600 n2643 n2644 n2623 VDD GND NOR2_X1
xU10601 n2625 n2626 n2624 VDD GND NOR2_X1
xU10602 n8363 n520 n2644 VDD GND NOR2_X1
xU10603 n2971 n2972 n7906 VDD GND NAND2_X1
xU10604 n2989 n2990 n2971 VDD GND NOR2_X1
xU10605 n2973 n2974 n2972 VDD GND NOR2_X1
xU10606 n8365 n490 n2990 VDD GND NOR2_X1
xU10607 n1135 n1136 n7852 VDD GND NAND2_X1
xU10608 n1156 n1157 n1135 VDD GND NOR2_X1
xU10609 n1137 n1138 n1136 VDD GND NOR2_X1
xU10610 n669 n8358 n1157 VDD GND NOR2_X1
xU10611 n1303 n1304 n7859 VDD GND NAND2_X1
xU10612 n1325 n1326 n1303 VDD GND NOR2_X1
xU10613 n1305 n1306 n1304 VDD GND NOR2_X1
xU10614 n8361 n650 n1326 VDD GND NOR2_X1
xU10615 n2547 n2548 n7891 VDD GND NAND2_X1
xU10616 n2570 n2571 n2547 VDD GND NOR2_X1
xU10617 n2549 n2550 n2548 VDD GND NOR2_X1
xU10618 n541 n8359 n2571 VDD GND NOR2_X1
xU10619 n2524 n2525 n7890 VDD GND NAND2_X1
xU10620 n2544 n2545 n2524 VDD GND NOR2_X1
xU10621 n2526 n2527 n2525 VDD GND NOR2_X1
xU10622 n542 n8360 n2545 VDD GND NOR2_X1
xU10623 n2776 n2777 n7900 VDD GND NAND2_X1
xU10624 n2800 n2801 n2776 VDD GND NOR2_X1
xU10625 n2778 n2779 n2777 VDD GND NOR2_X1
xU10626 n8364 n513 n2801 VDD GND NOR2_X1
xU10627 n1159 n1160 n7853 VDD GND NAND2_X1
xU10628 n1176 n1177 n1159 VDD GND NOR2_X1
xU10629 n1161 n1162 n1160 VDD GND NOR2_X1
xU10630 n668 n8358 n1177 VDD GND NOR2_X1
xU10631 n2727 n2728 n7898 VDD GND NAND2_X1
xU10632 n2749 n2750 n2727 VDD GND NOR2_X1
xU10633 n2729 n2730 n2728 VDD GND NOR2_X1
xU10634 n8364 n516 n2750 VDD GND NOR2_X1
xU10635 n1744 n1745 n7875 VDD GND NAND2_X1
xU10636 n1805 n1806 n1744 VDD GND NOR2_X1
xU10637 n1746 n1747 n1745 VDD GND NOR2_X1
xU10638 n8362 n594 n1806 VDD GND NOR2_X1
xU10639 n2404 n2405 n7885 VDD GND NAND2_X1
xU10640 n2427 n2428 n2404 VDD GND NOR2_X1
xU10641 n2406 n2407 n2405 VDD GND NOR2_X1
xU10642 n8363 n561 n2428 VDD GND NOR2_X1
xU10643 n1443 n1444 n7865 VDD GND NAND2_X1
xU10644 n1470 n1471 n1443 VDD GND NOR2_X1
xU10645 n1445 n1446 n1444 VDD GND NOR2_X1
xU10646 n8362 n625 n1471 VDD GND NOR2_X1
xU10647 n1496 n1497 n7867 VDD GND NAND2_X1
xU10648 n1522 n1523 n1496 VDD GND NOR2_X1
xU10649 n1498 n1499 n1497 VDD GND NOR2_X1
xU10650 n8363 n621 n1523 VDD GND NOR2_X1
xU10651 n1525 n1526 n7868 VDD GND NAND2_X1
xU10652 n1550 n1551 n1525 VDD GND NOR2_X1
xU10653 n1527 n1528 n1526 VDD GND NOR2_X1
xU10654 n8361 n618 n1551 VDD GND NOR2_X1
xU10655 n2899 n2900 n7905 VDD GND NAND2_X1
xU10656 n2968 n2969 n2899 VDD GND NOR2_X1
xU10657 n2901 n2902 n2900 VDD GND NOR2_X1
xU10658 n8365 n492 n2969 VDD GND NOR2_X1
xU10659 n2992 n2993 n7907 VDD GND NAND2_X1
xU10660 n3051 n3052 n2992 VDD GND NOR2_X1
xU10661 n2994 n2995 n2993 VDD GND NOR2_X1
xU10662 n8365 n489 n3052 VDD GND NOR2_X1
xU10663 n2290 n2291 n7881 VDD GND NAND2_X1
xU10664 n2315 n2316 n2290 VDD GND NOR2_X1
xU10665 n2292 n2293 n2291 VDD GND NOR2_X1
xU10666 n8363 n568 n2316 VDD GND NOR2_X1
xU10667 n2373 n2374 n7884 VDD GND NAND2_X1
xU10668 n2401 n2402 n2373 VDD GND NOR2_X1
xU10669 n2375 n2376 n2374 VDD GND NOR2_X1
xU10670 n8363 n563 n2402 VDD GND NOR2_X1
xU10671 n5524 n5525 n7972 VDD GND NAND2_X1
xU10672 n5576 n5577 n5524 VDD GND NOR2_X1
xU10673 n5526 n5527 n5525 VDD GND NOR2_X1
xU10674 n190 n8357 n5577 VDD GND NOR2_X1
xU10675 n2646 n2647 n7895 VDD GND NAND2_X1
xU10676 n2667 n2668 n2646 VDD GND NOR2_X1
xU10677 n2648 n2649 n2647 VDD GND NOR2_X1
xU10678 n8364 n519 n2668 VDD GND NOR2_X1
xU10679 n1033 n1034 n7848 VDD GND NAND2_X1
xU10680 n1051 n1052 n1033 VDD GND NOR2_X1
xU10681 n1035 n1036 n1034 VDD GND NOR2_X1
xU10682 n678 n8358 n1052 VDD GND NOR2_X1
xU10683 n1054 n1055 n7849 VDD GND NAND2_X1
xU10684 n1079 n1080 n1054 VDD GND NOR2_X1
xU10685 n1056 n1057 n1055 VDD GND NOR2_X1
xU10686 n677 n8357 n1080 VDD GND NOR2_X1
xU10687 n2454 n2455 n7887 VDD GND NAND2_X1
xU10688 n2472 n2473 n2454 VDD GND NOR2_X1
xU10689 n2456 n2457 n2455 VDD GND NOR2_X1
xU10690 n545 n8359 n2473 VDD GND NOR2_X1
xU10691 n3663 n3664 n7918 VDD GND NAND2_X1
xU10692 n3683 n3684 n3663 VDD GND NOR2_X1
xU10693 n3665 n3666 n3664 VDD GND NOR2_X1
xU10694 n8366 n443 n3684 VDD GND NOR2_X1
xU10695 n3884 n3885 n7927 VDD GND NAND2_X1
xU10696 n3904 n3905 n3884 VDD GND NOR2_X1
xU10697 n3886 n3887 n3885 VDD GND NOR2_X1
xU10698 n417 n8359 n3905 VDD GND NOR2_X1
xU10699 n3464 n3465 n7910 VDD GND NAND2_X1
xU10700 n3487 n3488 n3464 VDD GND NOR2_X1
xU10701 n3466 n3467 n3465 VDD GND NOR2_X1
xU10702 n8365 n468 n3488 VDD GND NOR2_X1
xU10703 n3686 n3687 n7919 VDD GND NAND2_X1
xU10704 n3708 n3709 n3686 VDD GND NOR2_X1
xU10705 n3688 n3689 n3687 VDD GND NOR2_X1
xU10706 n8366 n442 n3709 VDD GND NOR2_X1
xU10707 n1421 n1422 n7864 VDD GND NAND2_X1
xU10708 n1440 n1441 n1421 VDD GND NOR2_X1
xU10709 n1423 n1424 n1422 VDD GND NOR2_X1
xU10710 n8361 n626 n1441 VDD GND NOR2_X1
xU10711 n3860 n3861 n7926 VDD GND NAND2_X1
xU10712 n3881 n3882 n3860 VDD GND NOR2_X1
xU10713 n3862 n3863 n3861 VDD GND NOR2_X1
xU10714 n418 n8360 n3882 VDD GND NOR2_X1
xU10715 n3641 n3642 n7917 VDD GND NAND2_X1
xU10716 n3660 n3661 n3641 VDD GND NOR2_X1
xU10717 n3643 n3644 n3642 VDD GND NOR2_X1
xU10718 n8366 n459 n3661 VDD GND NOR2_X1
xU10719 n3618 n3619 n7916 VDD GND NAND2_X1
xU10720 n3638 n3639 n3618 VDD GND NOR2_X1
xU10721 n3620 n3621 n3619 VDD GND NOR2_X1
xU10722 n8366 n460 n3639 VDD GND NOR2_X1
xU10723 n3515 n3516 n7912 VDD GND NAND2_X1
xU10724 n3534 n3535 n3515 VDD GND NOR2_X1
xU10725 n3517 n3518 n3516 VDD GND NOR2_X1
xU10726 n8365 n466 n3535 VDD GND NOR2_X1
xU10727 n3711 n3712 n7920 VDD GND NAND2_X1
xU10728 n3729 n3730 n3711 VDD GND NOR2_X1
xU10729 n3713 n3714 n3712 VDD GND NOR2_X1
xU10730 n8366 n441 n3730 VDD GND NOR2_X1
xU10731 n4083 n4084 n7935 VDD GND NAND2_X1
xU10732 n4107 n4108 n4083 VDD GND NOR2_X1
xU10733 n4085 n4086 n4084 VDD GND NOR2_X1
xU10734 n8367 n394 n4108 VDD GND NOR2_X1
xU10735 n2870 n2871 n7904 VDD GND NAND2_X1
xU10736 n2896 n2897 n2870 VDD GND NOR2_X1
xU10737 n2872 n2873 n2871 VDD GND NOR2_X1
xU10738 n8365 n493 n2897 VDD GND NOR2_X1
xU10739 n2266 n2267 n7880 VDD GND NAND2_X1
xU10740 n2287 n2288 n2266 VDD GND NOR2_X1
xU10741 n2268 n2269 n2267 VDD GND NOR2_X1
xU10742 n8362 n570 n2288 VDD GND NOR2_X1
xU10743 n3732 n3733 n7921 VDD GND NAND2_X1
xU10744 n3753 n3754 n3732 VDD GND NOR2_X1
xU10745 n3734 n3735 n3733 VDD GND NOR2_X1
xU10746 n8366 n440 n3754 VDD GND NOR2_X1
xU10747 n1205 n1206 n7855 VDD GND NAND2_X1
xU10748 n1226 n1227 n1205 VDD GND NOR2_X1
xU10749 n1207 n1208 n1206 VDD GND NOR2_X1
xU10750 n8362 n655 n1227 VDD GND NOR2_X1
xU10751 n4060 n4061 n7934 VDD GND NAND2_X1
xU10752 n4080 n4081 n4060 VDD GND NOR2_X1
xU10753 n4062 n4063 n4061 VDD GND NOR2_X1
xU10754 n8367 n395 n4081 VDD GND NOR2_X1
xU10755 n2241 n2242 n7879 VDD GND NAND2_X1
xU10756 n2263 n2264 n2241 VDD GND NOR2_X1
xU10757 n2243 n2244 n2242 VDD GND NOR2_X1
xU10758 n8363 n571 n2264 VDD GND NOR2_X1
xU10759 n3927 n3928 n7929 VDD GND NAND2_X1
xU10760 n3954 n3955 n3927 VDD GND NOR2_X1
xU10761 n3929 n3930 n3928 VDD GND NOR2_X1
xU10762 n415 n8359 n3955 VDD GND NOR2_X1
xU10763 n1374 n1375 n7862 VDD GND NAND2_X1
xU10764 n1395 n1396 n1374 VDD GND NOR2_X1
xU10765 n1376 n1377 n1375 VDD GND NOR2_X1
xU10766 n8361 n628 n1396 VDD GND NOR2_X1
xU10767 n2499 n2500 n7889 VDD GND NAND2_X1
xU10768 n2521 n2522 n2499 VDD GND NOR2_X1
xU10769 n2501 n2502 n2500 VDD GND NOR2_X1
xU10770 n543 n8359 n2522 VDD GND NOR2_X1
xU10771 n2430 n2431 n7886 VDD GND NAND2_X1
xU10772 n2451 n2452 n2430 VDD GND NOR2_X1
xU10773 n2432 n2433 n2431 VDD GND NOR2_X1
xU10774 n546 n8360 n2452 VDD GND NOR2_X1
xU10775 n1723 n1724 n7874 VDD GND NAND2_X1
xU10776 n1741 n1742 n1723 VDD GND NOR2_X1
xU10777 n1725 n1726 n1724 VDD GND NOR2_X1
xU10778 n8362 n595 n1742 VDD GND NOR2_X1
xU10779 n1328 n1329 n7860 VDD GND NAND2_X1
xU10780 n1352 n1353 n1328 VDD GND NOR2_X1
xU10781 n1330 n1331 n1329 VDD GND NOR2_X1
xU10782 n8361 n647 n1353 VDD GND NOR2_X1
xU10783 n2670 n2671 n7896 VDD GND NAND2_X1
xU10784 n2693 n2694 n2670 VDD GND NOR2_X1
xU10785 n2672 n2673 n2671 VDD GND NOR2_X1
xU10786 n8364 n518 n2694 VDD GND NOR2_X1
xU10787 n2752 n2753 n7899 VDD GND NAND2_X1
xU10788 n2773 n2774 n2752 VDD GND NOR2_X1
xU10789 n2754 n2755 n2753 VDD GND NOR2_X1
xU10790 n8364 n515 n2774 VDD GND NOR2_X1
xU10791 n2803 n2804 n7901 VDD GND NAND2_X1
xU10792 n2820 n2821 n2803 VDD GND NOR2_X1
xU10793 n2805 n2806 n2804 VDD GND NOR2_X1
xU10794 n8364 n511 n2821 VDD GND NOR2_X1
xU10795 n2345 n2346 n7883 VDD GND NAND2_X1
xU10796 n2370 n2371 n2345 VDD GND NOR2_X1
xU10797 n2347 n2348 n2346 VDD GND NOR2_X1
xU10798 n8363 n565 n2371 VDD GND NOR2_X1
xU10799 n4110 n4111 n7936 VDD GND NAND2_X1
xU10800 n4137 n4138 n4110 VDD GND NOR2_X1
xU10801 n4112 n4113 n4111 VDD GND NOR2_X1
xU10802 n8367 n393 n4138 VDD GND NOR2_X1
xU10803 n3537 n3538 n7913 VDD GND NAND2_X1
xU10804 n3560 n3561 n3537 VDD GND NOR2_X1
xU10805 n3539 n3540 n3538 VDD GND NOR2_X1
xU10806 n8365 n465 n3561 VDD GND NOR2_X1
xU10807 n3490 n3491 n7911 VDD GND NAND2_X1
xU10808 n3512 n3513 n3490 VDD GND NOR2_X1
xU10809 n3492 n3493 n3491 VDD GND NOR2_X1
xU10810 n8365 n467 n3513 VDD GND NOR2_X1
xU10811 n4140 n4141 n7937 VDD GND NAND2_X1
xU10812 n4210 n4211 n4140 VDD GND NOR2_X1
xU10813 n4142 n4143 n4141 VDD GND NOR2_X1
xU10814 n8367 n392 n4211 VDD GND NOR2_X1
xU10815 n3054 n3055 n7908 VDD GND NAND2_X1
xU10816 n3106 n3107 n3054 VDD GND NOR2_X1
xU10817 n3056 n3057 n3055 VDD GND NOR2_X1
xU10818 n8365 n485 n3107 VDD GND NOR2_X1
xU10819 n1575 n1576 n7870 VDD GND NAND2_X1
xU10820 n1594 n1595 n1575 VDD GND NOR2_X1
xU10821 n1577 n1578 n1576 VDD GND NOR2_X1
xU10822 n8361 n600 n1595 VDD GND NOR2_X1
xU10823 n4234 n4235 n7939 VDD GND NAND2_X1
xU10824 n4295 n4296 n4234 VDD GND NOR2_X1
xU10825 n4236 n4237 n4235 VDD GND NOR2_X1
xU10826 n8367 n389 n4296 VDD GND NOR2_X1
xU10827 n2845 n2846 n7903 VDD GND NAND2_X1
xU10828 n2867 n2868 n2845 VDD GND NOR2_X1
xU10829 n2847 n2848 n2846 VDD GND NOR2_X1
xU10830 n8364 n494 n2868 VDD GND NOR2_X1
xU10831 n1652 n1653 n7873 VDD GND NAND2_X1
xU10832 n1720 n1721 n1652 VDD GND NOR2_X1
xU10833 n1654 n1655 n1653 VDD GND NOR2_X1
xU10834 n8363 n597 n1721 VDD GND NOR2_X1
xU10835 n4298 n4299 n7940 VDD GND NAND2_X1
xU10836 n4340 n4341 n4298 VDD GND NOR2_X1
xU10837 n4300 n4301 n4299 VDD GND NOR2_X1
xU10838 n8367 n388 n4341 VDD GND NOR2_X1
xU10839 n4039 n4040 n7933 VDD GND NAND2_X1
xU10840 n4057 n4058 n4039 VDD GND NOR2_X1
xU10841 n4041 n4042 n4040 VDD GND NOR2_X1
xU10842 n409 n8358 n4058 VDD GND NOR2_X1
xU10843 n3982 n3983 n7931 VDD GND NAND2_X1
xU10844 n4005 n4006 n3982 VDD GND NOR2_X1
xU10845 n3984 n3985 n3983 VDD GND NOR2_X1
xU10846 n412 n8358 n4006 VDD GND NOR2_X1
xU10847 n3590 n3591 n7915 VDD GND NAND2_X1
xU10848 n3615 n3616 n3590 VDD GND NOR2_X1
xU10849 n3592 n3593 n3591 VDD GND NOR2_X1
xU10850 n8366 n462 n3616 VDD GND NOR2_X1
xU10851 n3907 n3908 n7928 VDD GND NAND2_X1
xU10852 n3924 n3925 n3907 VDD GND NOR2_X1
xU10853 n3909 n3910 n3908 VDD GND NOR2_X1
xU10854 n416 n8360 n3925 VDD GND NOR2_X1
xU10855 n4008 n4009 n7932 VDD GND NAND2_X1
xU10856 n4036 n4037 n4008 VDD GND NOR2_X1
xU10857 n4010 n4011 n4009 VDD GND NOR2_X1
xU10858 n411 n8359 n4037 VDD GND NOR2_X1
xU10859 n3563 n3564 n7914 VDD GND NAND2_X1
xU10860 n3587 n3588 n3563 VDD GND NOR2_X1
xU10861 n3565 n3566 n3564 VDD GND NOR2_X1
xU10862 n8366 n463 n3588 VDD GND NOR2_X1
xU10863 n982 n983 n7846 VDD GND NAND2_X1
xU10864 n1005 n1006 n982 VDD GND NOR2_X1
xU10865 n984 n985 n983 VDD GND NOR2_X1
xU10866 n680 n8359 n1006 VDD GND NOR2_X1
xU10867 n4343 n4344 n7941 VDD GND NAND2_X1
xU10868 n4696 n4697 n4343 VDD GND NOR2_X1
xU10869 n4345 n4346 n4344 VDD GND NOR2_X1
xU10870 n8367 n386 n4697 VDD GND NOR2_X1
xU10871 n2318 n2319 n7882 VDD GND NAND2_X1
xU10872 n2342 n2343 n2318 VDD GND NOR2_X1
xU10873 n2320 n2321 n2319 VDD GND NOR2_X1
xU10874 n8363 n566 n2343 VDD GND NOR2_X1
xU10875 n3812 n3813 n7924 VDD GND NAND2_X1
xU10876 n3837 n3838 n3812 VDD GND NOR2_X1
xU10877 n3814 n3815 n3813 VDD GND NOR2_X1
xU10878 n8367 n434 n3838 VDD GND NOR2_X1
xU10879 n2573 n2574 n7892 VDD GND NAND2_X1
xU10880 n2598 n2599 n2573 VDD GND NOR2_X1
xU10881 n2575 n2576 n2574 VDD GND NOR2_X1
xU10882 n539 n8360 n2599 VDD GND NOR2_X1
xU10883 n3840 n3841 n7925 VDD GND NAND2_X1
xU10884 n3857 n3858 n3840 VDD GND NOR2_X1
xU10885 n3842 n3843 n3841 VDD GND NOR2_X1
xU10886 n8367 n433 n3858 VDD GND NOR2_X1
xU10887 n1276 n1277 n7858 VDD GND NAND2_X1
xU10888 n1300 n1301 n1276 VDD GND NOR2_X1
xU10889 n1278 n1279 n1277 VDD GND NOR2_X1
xU10890 n8360 n651 n1301 VDD GND NOR2_X1
xU10891 n2601 n2602 n7893 VDD GND NAND2_X1
xU10892 n2620 n2621 n2601 VDD GND NOR2_X1
xU10893 n2603 n2604 n2602 VDD GND NOR2_X1
xU10894 n538 n8359 n2621 VDD GND NOR2_X1
xU10895 n3756 n3757 n7922 VDD GND NAND2_X1
xU10896 n3778 n3779 n3756 VDD GND NOR2_X1
xU10897 n3758 n3759 n3757 VDD GND NOR2_X1
xU10898 n8366 n437 n3779 VDD GND NOR2_X1
xU10899 n3957 n3958 n7930 VDD GND NAND2_X1
xU10900 n3979 n3980 n3957 VDD GND NOR2_X1
xU10901 n3959 n3960 n3958 VDD GND NOR2_X1
xU10902 n413 n8359 n3980 VDD GND NOR2_X1
xU10903 n1473 n1474 n7866 VDD GND NAND2_X1
xU10904 n1493 n1494 n1473 VDD GND NOR2_X1
xU10905 n1475 n1476 n1474 VDD GND NOR2_X1
xU10906 n8361 n622 n1494 VDD GND NOR2_X1
xU10907 n4213 n4214 n7938 VDD GND NAND2_X1
xU10908 n4231 n4232 n4213 VDD GND NOR2_X1
xU10909 n4215 n4216 n4214 VDD GND NOR2_X1
xU10910 n8367 n390 n4232 VDD GND NOR2_X1
xU10911 n3109 n3110 n7909 VDD GND NAND2_X1
xU10912 n3461 n3462 n3109 VDD GND NOR2_X1
xU10913 n3111 n3112 n3110 VDD GND NOR2_X1
xU10914 n8365 n483 n3462 VDD GND NOR2_X1
xU10915 n2650 n931 n2649 VDD GND NOR2_X1
xU10916 n2651 n2652 n2650 VDD GND NOR2_X1
xU10917 n227 n8411 n2652 VDD GND NOR2_X1
xU10918 n218 n8378 n2651 VDD GND NOR2_X1
xU10919 n1402 n963 n1401 VDD GND NOR2_X1
xU10920 n1403 n1404 n1402 VDD GND NOR2_X1
xU10921 n1405 n8406 n1404 VDD GND NOR2_X1
xU10922 n180 n8384 n1403 VDD GND NOR2_X1
xU10923 \AES_Comp_ENCa/KrgX_124 n1063 n1056 VDD GND NOR2_X1
xU10924 n1064 n1065 n1063 VDD GND NOR2_X1
xU10925 n662 n8402 n1065 VDD GND NOR2_X1
xU10926 n168 n8387 n1064 VDD GND NOR2_X1
xU10927 \AES_Comp_ENCa/KrgX_55 n3672 n3665 VDD GND NOR2_X1
xU10928 n3673 n3674 n3672 VDD GND NOR2_X1
xU10929 n3670 n8408 n3674 VDD GND NOR2_X1
xU10930 n295 n8381 n3673 VDD GND NOR2_X1
xU10931 \AES_Comp_ENCa/KrgX_63 n3473 n3466 VDD GND NOR2_X1
xU10932 n3474 n3475 n3473 VDD GND NOR2_X1
xU10933 n3471 n8410 n3475 VDD GND NOR2_X1
xU10934 n286 n8380 n3474 VDD GND NOR2_X1
xU10935 \AES_Comp_ENCa/KrgX_23 n4908 n4901 VDD GND NOR2_X1
xU10936 n4909 n4910 n4908 VDD GND NOR2_X1
xU10937 n4906 n8404 n4910 VDD GND NOR2_X1
xU10938 n327 n8385 n4909 VDD GND NOR2_X1
xU10939 n3622 n910 n3621 VDD GND NOR2_X1
xU10940 n3623 n3624 n3622 VDD GND NOR2_X1
xU10941 n3625 n8409 n3624 VDD GND NOR2_X1
xU10942 n266 n8381 n3623 VDD GND NOR2_X1
xU10943 \AES_Comp_ENCa/KrgX_71 n2832 n2825 VDD GND NOR2_X1
xU10944 n2833 n2834 n2832 VDD GND NOR2_X1
xU10945 n2830 n8410 n2834 VDD GND NOR2_X1
xU10946 n208 n8379 n2833 VDD GND NOR2_X1
xU10947 n4087 n891 n4086 VDD GND NOR2_X1
xU10948 n4088 n4089 n4087 VDD GND NOR2_X1
xU10949 n475 n8406 n4089 VDD GND NOR2_X1
xU10950 n292 n8383 n4088 VDD GND NOR2_X1
xU10951 n1209 n971 n1208 VDD GND NOR2_X1
xU10952 n1210 n1211 n1209 VDD GND NOR2_X1
xU10953 n531 n8404 n1211 VDD GND NOR2_X1
xU10954 n174 n8386 n1210 VDD GND NOR2_X1
xU10955 \AES_Comp_ENCa/KrgX_67 n2980 n2973 VDD GND NOR2_X1
xU10956 n2981 n2982 n2980 VDD GND NOR2_X1
xU10957 n580 n8410 n2982 VDD GND NOR2_X1
xU10958 n204 n8380 n2981 VDD GND NOR2_X1
xU10959 \AES_Comp_ENCa/KrgX_123 n1091 n1084 VDD GND NOR2_X1
xU10960 n1092 n1093 n1091 VDD GND NOR2_X1
xU10961 n664 n8403 n1093 VDD GND NOR2_X1
xU10962 n178 n8387 n1092 VDD GND NOR2_X1
xU10963 n1139 n974 n1138 VDD GND NOR2_X1
xU10964 n1140 n1141 n1139 VDD GND NOR2_X1
xU10965 n660 n8403 n1141 VDD GND NOR2_X1
xU10966 n156 n8387 n1140 VDD GND NOR2_X1
xU10967 \AES_Comp_ENCa/KrgX_87 n2439 n2432 VDD GND NOR2_X1
xU10968 n2440 n2441 n2439 VDD GND NOR2_X1
xU10969 n2437 n8412 n2441 VDD GND NOR2_X1
xU10970 n212 n8378 n2440 VDD GND NOR2_X1
xU10971 \AES_Comp_ENCa/KrgX_83 n2532 n2526 VDD GND NOR2_X1
xU10972 n2533 n2534 n2532 VDD GND NOR2_X1
xU10973 n2283 n8412 n2534 VDD GND NOR2_X1
xU10974 n214 n8378 n2533 VDD GND NOR2_X1
xU10975 \AES_Comp_ENCa/KrgX_12 n5166 n5159 VDD GND NOR2_X1
xU10976 n5167 n5168 n5166 VDD GND NOR2_X1
xU10977 n5164 n8403 n5168 VDD GND NOR2_X1
xU10978 n333 n8386 n5167 VDD GND NOR2_X1
xU10979 n5240 n840 n5239 VDD GND NOR2_X1
xU10980 n5241 n5242 n5240 VDD GND NOR2_X1
xU10981 n500 n8403 n5242 VDD GND NOR2_X1
xU10982 n317 n8387 n5241 VDD GND NOR2_X1
xU10983 \AES_Comp_ENCa/KrgX_90 n2354 n2347 VDD GND NOR2_X1
xU10984 n2355 n2356 n2354 VDD GND NOR2_X1
xU10985 n2352 n8411 n2356 VDD GND NOR2_X1
xU10986 n207 n8379 n2355 VDD GND NOR2_X1
xU10987 n1601 n955 n1600 VDD GND NOR2_X1
xU10988 n1602 n1603 n1601 VDD GND NOR2_X1
xU10989 n173 n8408 n1603 VDD GND NOR2_X1
xU10990 n162 n8382 n1602 VDD GND NOR2_X1
xU10991 \AES_Comp_ENCa/KrgX_27 n4808 n4802 VDD GND NOR2_X1
xU10992 n4809 n4810 n4808 VDD GND NOR2_X1
xU10993 n4811 n8405 n4810 VDD GND NOR2_X1
xU10994 n348 n8385 n4809 VDD GND NOR2_X1
xU10995 \AES_Comp_ENCa/KrgX_122 n1116 n1109 VDD GND NOR2_X1
xU10996 n1117 n1118 n1116 VDD GND NOR2_X1
xU10997 n657 n8403 n1118 VDD GND NOR2_X1
xU10998 n150 n8387 n1117 VDD GND NOR2_X1
xU10999 n2479 n938 n2478 VDD GND NOR2_X1
xU11000 n2480 n2481 n2479 VDD GND NOR2_X1
xU11001 n2482 n8410 n2481 VDD GND NOR2_X1
xU11002 n201 n8383 n2480 VDD GND NOR2_X1
xU11003 \AES_Comp_ENCa/KrgX_75 n2735 n2729 VDD GND NOR2_X1
xU11004 n2736 n2737 n2735 VDD GND NOR2_X1
xU11005 n2738 n8411 n2737 VDD GND NOR2_X1
xU11006 n225 n8379 n2736 VDD GND NOR2_X1
xU11007 \AES_Comp_ENCa/KrgX_34 n4243 n4236 VDD GND NOR2_X1
xU11008 n4244 n4245 n4243 VDD GND NOR2_X1
xU11009 n4241 n8406 n4245 VDD GND NOR2_X1
xU11010 n4242 n8384 n4244 VDD GND NOR2_X1
xU11011 n2849 n923 n2848 VDD GND NOR2_X1
xU11012 n2850 n2851 n2849 VDD GND NOR2_X1
xU11013 n2261 n8410 n2851 VDD GND NOR2_X1
xU11014 n223 n8379 n2850 VDD GND NOR2_X1
xU11015 n5528 n825 n5527 VDD GND NOR2_X1
xU11016 n5529 n5530 n5528 VDD GND NOR2_X1
xU11017 n5057 n8402 n5530 VDD GND NOR2_X1
xU11018 n337 n8387 n5529 VDD GND NOR2_X1
xU11019 n4858 n876 n4857 VDD GND NOR2_X1
xU11020 n4859 n4860 n4858 VDD GND NOR2_X1
xU11021 n4861 n8405 n4860 VDD GND NOR2_X1
xU11022 n314 n8385 n4859 VDD GND NOR2_X1
xU11023 n4302 n886 n4301 VDD GND NOR2_X1
xU11024 n4303 n4304 n4302 VDD GND NOR2_X1
xU11025 n3637 n8406 n4304 VDD GND NOR2_X1
xU11026 n274 n8384 n4303 VDD GND NOR2_X1
xU11027 \AES_Comp_ENCa/KrgX_106 n1505 n1498 VDD GND NOR2_X1
xU11028 n1506 n1507 n1505 VDD GND NOR2_X1
xU11029 n1503 n8407 n1507 VDD GND NOR2_X1
xU11030 n142 n8383 n1506 VDD GND NOR2_X1
xU11031 \AES_Comp_ENCa/KrgX_58 n3599 n3592 VDD GND NOR2_X1
xU11032 n3600 n3601 n3599 VDD GND NOR2_X1
xU11033 n3597 n8409 n3601 VDD GND NOR2_X1
xU11034 n294 n8381 n3600 VDD GND NOR2_X1
xU11035 n4012 n894 n4011 VDD GND NOR2_X1
xU11036 n4013 n4014 n4012 VDD GND NOR2_X1
xU11037 n4015 n8407 n4014 VDD GND NOR2_X1
xU11038 n275 n8383 n4013 VDD GND NOR2_X1
xU11039 \AES_Comp_ENCa/KrgX_7 n5298 n5291 VDD GND NOR2_X1
xU11040 n5299 n5300 n5298 VDD GND NOR2_X1
xU11041 n5296 n8402 n5300 VDD GND NOR2_X1
xU11042 n316 n8386 n5299 VDD GND NOR2_X1
xU11043 \AES_Comp_ENCa/KrgX_91 n2327 n2320 VDD GND NOR2_X1
xU11044 n2328 n2329 n2327 VDD GND NOR2_X1
xU11045 n2325 n8411 n2329 VDD GND NOR2_X1
xU11046 n202 n8379 n2328 VDD GND NOR2_X1
xU11047 n2377 n942 n2376 VDD GND NOR2_X1
xU11048 n2378 n2379 n2377 VDD GND NOR2_X1
xU11049 n550 n8411 n2379 VDD GND NOR2_X1
xU11050 n236 n8378 n2378 VDD GND NOR2_X1
xU11051 n3844 n901 n3843 VDD GND NOR2_X1
xU11052 n3845 n3846 n3844 VDD GND NOR2_X1
xU11053 n3847 n8408 n3846 VDD GND NOR2_X1
xU11054 n279 n8382 n3845 VDD GND NOR2_X1
xU11055 n5046 n857 n5045 VDD GND NOR2_X1
xU11056 n5047 n5048 n5046 VDD GND NOR2_X1
xU11057 n632 n8404 n5048 VDD GND NOR2_X1
xU11058 n318 n8386 n5047 VDD GND NOR2_X1
xU11059 n2605 n933 n2604 VDD GND NOR2_X1
xU11060 n2606 n2607 n2605 VDD GND NOR2_X1
xU11061 n2608 n8412 n2607 VDD GND NOR2_X1
xU11062 n222 n8378 n2606 VDD GND NOR2_X1
xU11063 \AES_Comp_ENCa/KrgX_35 n4221 n4215 VDD GND NOR2_X1
xU11064 n4222 n4223 n4221 VDD GND NOR2_X1
xU11065 n478 n8406 n4223 VDD GND NOR2_X1
xU11066 n259 n8384 n4222 VDD GND NOR2_X1
xU11067 \AES_Comp_ENCa/KrgX_127 n993 n984 VDD GND NOR2_X1
xU11068 n994 n995 n993 VDD GND NOR2_X1
xU11069 n658 n8402 n995 VDD GND NOR2_X1
xU11070 n151 n8388 n994 VDD GND NOR2_X1
xU11071 \AES_Comp_ENCa/KrgX_3 n5445 n5439 VDD GND NOR2_X1
xU11072 n5446 n5447 n5445 VDD GND NOR2_X1
xU11073 n372 n8402 n5447 VDD GND NOR2_X1
xU11074 n338 n8388 n5446 VDD GND NOR2_X1
xU11075 n4238 n887 n4237 VDD GND NOR2_X1
xU11076 n4239 n4240 n4238 VDD GND NOR2_X1
xU11077 n8430 n476 n4240 VDD GND NOR2_X1
xU11078 n8395 n282 n4239 VDD GND NOR2_X1
xU11079 \AES_Comp_ENCa/KrgX_101 n1630 n1624 VDD GND NOR2_X1
xU11080 n1631 n1632 n1630 VDD GND NOR2_X1
xU11081 n8425 n1612 n1632 VDD GND NOR2_X1
xU11082 n8390 n167 n1631 VDD GND NOR2_X1
xU11083 \AES_Comp_ENCa/KrgX_125 n1042 n1035 VDD GND NOR2_X1
xU11084 n1043 n1044 n1042 VDD GND NOR2_X1
xU11085 n8426 n661 n1044 VDD GND NOR2_X1
xU11086 n8391 n160 n1043 VDD GND NOR2_X1
xU11087 \AES_Comp_ENCa/KrgX_86 n2463 n2456 VDD GND NOR2_X1
xU11088 n2464 n2465 n2463 VDD GND NOR2_X1
xU11089 n8426 n425 n2465 VDD GND NOR2_X1
xU11090 n8391 n219 n2464 VDD GND NOR2_X1
xU11091 n2221 n948 n2220 VDD GND NOR2_X1
xU11092 n2222 n2223 n2221 VDD GND NOR2_X1
xU11093 n8424 n551 n2223 VDD GND NOR2_X1
xU11094 n8390 n213 n2222 VDD GND NOR2_X1
xU11095 \AES_Comp_ENCa/KrgX_46 n3892 n3886 VDD GND NOR2_X1
xU11096 n3893 n3894 n3892 VDD GND NOR2_X1
xU11097 n8429 n3895 n3894 VDD GND NOR2_X1
xU11098 n8395 n293 n3893 VDD GND NOR2_X1
xU11099 n2627 n932 n2626 VDD GND NOR2_X1
xU11100 n2628 n2629 n2627 VDD GND NOR2_X1
xU11101 n8427 n209 n2629 VDD GND NOR2_X1
xU11102 n8392 n226 n2628 VDD GND NOR2_X1
xU11103 \AES_Comp_ENCa/KrgX_54 n3695 n3688 VDD GND NOR2_X1
xU11104 n3696 n3697 n3695 VDD GND NOR2_X1
xU11105 n8429 n296 n3697 VDD GND NOR2_X1
xU11106 n8394 n271 n3696 VDD GND NOR2_X1
xU11107 \AES_Comp_ENCa/KrgX_109 n1430 n1423 VDD GND NOR2_X1
xU11108 n1431 n1432 n1430 VDD GND NOR2_X1
xU11109 n8423 n398 n1432 VDD GND NOR2_X1
xU11110 n8388 n176 n1431 VDD GND NOR2_X1
xU11111 n3864 n900 n3863 VDD GND NOR2_X1
xU11112 n3865 n3866 n3864 VDD GND NOR2_X1
xU11113 n8429 n3867 n3866 VDD GND NOR2_X1
xU11114 n8394 n280 n3865 VDD GND NOR2_X1
xU11115 \AES_Comp_ENCa/KrgX_56 n3650 n3643 VDD GND NOR2_X1
xU11116 n3651 n3652 n3650 VDD GND NOR2_X1
xU11117 n8428 n451 n3652 VDD GND NOR2_X1
xU11118 n8394 n264 n3651 VDD GND NOR2_X1
xU11119 \AES_Comp_ENCa/KrgX_61 n3523 n3517 VDD GND NOR2_X1
xU11120 n3524 n3525 n3523 VDD GND NOR2_X1
xU11121 n8428 n447 n3525 VDD GND NOR2_X1
xU11122 n8393 n261 n3524 VDD GND NOR2_X1
xU11123 \AES_Comp_ENCa/KrgX_53 n3719 n3713 VDD GND NOR2_X1
xU11124 n3720 n3721 n3719 VDD GND NOR2_X1
xU11125 n8429 n3701 n3721 VDD GND NOR2_X1
xU11126 n8394 n289 n3720 VDD GND NOR2_X1
xU11127 \AES_Comp_ENCa/KrgX_22 n4932 n4925 VDD GND NOR2_X1
xU11128 n4933 n4934 n4932 VDD GND NOR2_X1
xU11129 n8431 n4930 n4934 VDD GND NOR2_X1
xU11130 n8396 n350 n4933 VDD GND NOR2_X1
xU11131 \AES_Comp_ENCa/KrgX_29 n4762 n4756 VDD GND NOR2_X1
xU11132 n4763 n4764 n4762 VDD GND NOR2_X1
xU11133 n8430 n323 n4764 VDD GND NOR2_X1
xU11134 n8396 n336 n4763 VDD GND NOR2_X1
xU11135 \AES_Comp_ENCa/KrgX_69 n2879 n2872 VDD GND NOR2_X1
xU11136 n2880 n2881 n2879 VDD GND NOR2_X1
xU11137 n8427 n574 n2881 VDD GND NOR2_X1
xU11138 n8393 n215 n2880 VDD GND NOR2_X1
xU11139 \AES_Comp_ENCa/KrgX_93 n2274 n2268 VDD GND NOR2_X1
xU11140 n2275 n2276 n2274 VDD GND NOR2_X1
xU11141 n8424 n2258 n2276 VDD GND NOR2_X1
xU11142 n8390 n216 n2275 VDD GND NOR2_X1
xU11143 n3736 n905 n3735 VDD GND NOR2_X1
xU11144 n3737 n3738 n3736 VDD GND NOR2_X1
xU11145 n8429 n3739 n3738 VDD GND NOR2_X1
xU11146 n8394 n265 n3737 VDD GND NOR2_X1
xU11147 n4973 n864 n4972 VDD GND NOR2_X1
xU11148 n4974 n4975 n4973 VDD GND NOR2_X1
xU11149 n8431 n4976 n4975 VDD GND NOR2_X1
xU11150 n8397 n334 n4974 VDD GND NOR2_X1
xU11151 \AES_Comp_ENCa/KrgX_30 n4738 n4731 VDD GND NOR2_X1
xU11152 n4739 n4740 n4738 VDD GND NOR2_X1
xU11153 n8430 n351 n4740 VDD GND NOR2_X1
xU11154 n8396 n324 n4739 VDD GND NOR2_X1
xU11155 n4064 n892 n4063 VDD GND NOR2_X1
xU11156 n4065 n4066 n4064 VDD GND NOR2_X1
xU11157 n8430 n3479 n4066 VDD GND NOR2_X1
xU11158 n8395 n278 n4065 VDD GND NOR2_X1
xU11159 \AES_Comp_ENCa/KrgX_94 n2250 n2243 VDD GND NOR2_X1
xU11160 n2251 n2252 n2250 VDD GND NOR2_X1
xU11161 n8424 n555 n2252 VDD GND NOR2_X1
xU11162 n8390 n224 n2251 VDD GND NOR2_X1
xU11163 n5215 n841 n5214 VDD GND NOR2_X1
xU11164 n5216 n5217 n5215 VDD GND NOR2_X1
xU11165 n8432 n502 n5217 VDD GND NOR2_X1
xU11166 n8397 n330 n5216 VDD GND NOR2_X1
xU11167 n1183 n972 n1182 VDD GND NOR2_X1
xU11168 n1184 n1185 n1183 VDD GND NOR2_X1
xU11169 n8426 n526 n1185 VDD GND NOR2_X1
xU11170 n8390 n147 n1184 VDD GND NOR2_X1
xU11171 n3931 n897 n3930 VDD GND NOR2_X1
xU11172 n3932 n3933 n3931 VDD GND NOR2_X1
xU11173 n8429 n3557 n3933 VDD GND NOR2_X1
xU11174 n8395 n288 n3932 VDD GND NOR2_X1
xU11175 n1378 n964 n1377 VDD GND NOR2_X1
xU11176 n1379 n1380 n1378 VDD GND NOR2_X1
xU11177 n8423 n400 n1380 VDD GND NOR2_X1
xU11178 n8389 n152 n1379 VDD GND NOR2_X1
xU11179 \AES_Comp_ENCa/KrgX_126 n1018 n1012 VDD GND NOR2_X1
xU11180 n1019 n1020 n1018 VDD GND NOR2_X1
xU11181 n8426 n1021 n1020 VDD GND NOR2_X1
xU11182 n8391 n175 n1019 VDD GND NOR2_X1
xU11183 n2503 n937 n2502 VDD GND NOR2_X1
xU11184 n2504 n2505 n2503 VDD GND NOR2_X1
xU11185 n8426 n420 n2505 VDD GND NOR2_X1
xU11186 n8392 n238 n2504 VDD GND NOR2_X1
xU11187 n5094 n847 n5093 VDD GND NOR2_X1
xU11188 n5095 n5096 n5094 VDD GND NOR2_X1
xU11189 n8432 n5097 n5096 VDD GND NOR2_X1
xU11190 n8397 n325 n5095 VDD GND NOR2_X1
xU11191 n1254 n969 n1253 VDD GND NOR2_X1
xU11192 n1255 n1256 n1254 VDD GND NOR2_X1
xU11193 n8425 n1257 n1256 VDD GND NOR2_X1
xU11194 n8389 n165 n1255 VDD GND NOR2_X1
xU11195 n1727 n952 n1726 VDD GND NOR2_X1
xU11196 n1728 n1729 n1727 VDD GND NOR2_X1
xU11197 n8424 n179 n1729 VDD GND NOR2_X1
xU11198 n8389 n163 n1728 VDD GND NOR2_X1
xU11199 n1307 n967 n1306 VDD GND NOR2_X1
xU11200 n1308 n1309 n1307 VDD GND NOR2_X1
xU11201 n8424 n1310 n1309 VDD GND NOR2_X1
xU11202 n8389 n146 n1308 VDD GND NOR2_X1
xU11203 n2551 n935 n2550 VDD GND NOR2_X1
xU11204 n2552 n2553 n2551 VDD GND NOR2_X1
xU11205 n8426 n2554 n2553 VDD GND NOR2_X1
xU11206 n8392 n211 n2552 VDD GND NOR2_X1
xU11207 n3785 n903 n3784 VDD GND NOR2_X1
xU11208 n3786 n3787 n3785 VDD GND NOR2_X1
xU11209 n8429 n3788 n3787 VDD GND NOR2_X1
xU11210 n8394 n276 n3786 VDD GND NOR2_X1
xU11211 \AES_Comp_ENCa/KrgX_21 n4954 n4948 VDD GND NOR2_X1
xU11212 n4955 n4956 n4954 VDD GND NOR2_X1
xU11213 n8431 n4957 n4956 VDD GND NOR2_X1
xU11214 n8396 n322 n4955 VDD GND NOR2_X1
xU11215 \AES_Comp_ENCa/KrgX_113 n1337 n1330 VDD GND NOR2_X1
xU11216 n1338 n1339 n1337 VDD GND NOR2_X1
xU11217 n8425 n524 n1339 VDD GND NOR2_X1
xU11218 n8389 n157 n1338 VDD GND NOR2_X1
xU11219 \AES_Comp_ENCa/KrgX_77 n2679 n2672 VDD GND NOR2_X1
xU11220 n2680 n2681 n2679 VDD GND NOR2_X1
xU11221 n8427 n2677 n2681 VDD GND NOR2_X1
xU11222 n8392 n230 n2680 VDD GND NOR2_X1
xU11223 \AES_Comp_ENCa/KrgX_14 n5122 n5115 VDD GND NOR2_X1
xU11224 n5123 n5124 n5122 VDD GND NOR2_X1
xU11225 n8432 n505 n5124 VDD GND NOR2_X1
xU11226 n8397 n349 n5123 VDD GND NOR2_X1
xU11227 n2756 n927 n2755 VDD GND NOR2_X1
xU11228 n2757 n2758 n2756 VDD GND NOR2_X1
xU11229 n8427 n2759 n2758 VDD GND NOR2_X1
xU11230 n8392 n235 n2757 VDD GND NOR2_X1
xU11231 \AES_Comp_ENCa/KrgX_8 n5275 n5268 VDD GND NOR2_X1
xU11232 n5276 n5277 n5275 VDD GND NOR2_X1
xU11233 n8432 n496 n5277 VDD GND NOR2_X1
xU11234 n8397 n340 n5276 VDD GND NOR2_X1
xU11235 \AES_Comp_ENCa/KrgX_73 n2785 n2778 VDD GND NOR2_X1
xU11236 n2786 n2787 n2785 VDD GND NOR2_X1
xU11237 n8427 n2783 n2787 VDD GND NOR2_X1
xU11238 n8392 n221 n2786 VDD GND NOR2_X1
xU11239 \AES_Comp_ENCa/KrgX_13 n5145 n5139 VDD GND NOR2_X1
xU11240 n5146 n5147 n5145 VDD GND NOR2_X1
xU11241 n8432 n5128 n5147 VDD GND NOR2_X1
xU11242 n8397 n321 n5146 VDD GND NOR2_X1
xU11243 n2700 n929 n2699 VDD GND NOR2_X1
xU11244 n2701 n2702 n2700 VDD GND NOR2_X1
xU11245 n8427 n231 n2702 VDD GND NOR2_X1
xU11246 n8392 n228 n2701 VDD GND NOR2_X1
xU11247 \AES_Comp_ENCa/KrgX_72 n2811 n2805 VDD GND NOR2_X1
xU11248 n2812 n2813 n2811 VDD GND NOR2_X1
xU11249 n8427 n199 n2813 VDD GND NOR2_X1
xU11250 n8393 n210 n2812 VDD GND NOR2_X1
xU11251 n4830 n878 n4829 VDD GND NOR2_X1
xU11252 n4831 n4832 n4830 VDD GND NOR2_X1
xU11253 n8431 n4833 n4832 VDD GND NOR2_X1
xU11254 n8396 n319 n4831 VDD GND NOR2_X1
xU11255 n4779 n880 n4778 VDD GND NOR2_X1
xU11256 n4780 n4781 n4779 VDD GND NOR2_X1
xU11257 n8431 n335 n4781 VDD GND NOR2_X1
xU11258 n8396 n329 n4780 VDD GND NOR2_X1
xU11259 \AES_Comp_ENCa/KrgX_24 n4888 n4881 VDD GND NOR2_X1
xU11260 n4889 n4890 n4888 VDD GND NOR2_X1
xU11261 n8431 n342 n4890 VDD GND NOR2_X1
xU11262 n8396 n326 n4889 VDD GND NOR2_X1
xU11263 \AES_Comp_ENCa/KrgX_37 n4118 n4112 VDD GND NOR2_X1
xU11264 n4119 n4120 n4118 VDD GND NOR2_X1
xU11265 n8430 n4098 n4120 VDD GND NOR2_X1
xU11266 n8395 n268 n4119 VDD GND NOR2_X1
xU11267 n3541 n913 n3540 VDD GND NOR2_X1
xU11268 n3542 n3543 n3541 VDD GND NOR2_X1
xU11269 n8428 n3530 n3543 VDD GND NOR2_X1
xU11270 n8393 n273 n3542 VDD GND NOR2_X1
xU11271 \AES_Comp_ENCa/KrgX_62 n3498 n3492 VDD GND NOR2_X1
xU11272 n3499 n3500 n3498 VDD GND NOR2_X1
xU11273 n8428 n3501 n3500 VDD GND NOR2_X1
xU11274 n8393 n272 n3499 VDD GND NOR2_X1
xU11275 n5022 n860 n5021 VDD GND NOR2_X1
xU11276 n5023 n5024 n5022 VDD GND NOR2_X1
xU11277 n8431 n634 n5024 VDD GND NOR2_X1
xU11278 n8397 n331 n5023 VDD GND NOR2_X1
xU11279 n4144 n889 n4143 VDD GND NOR2_X1
xU11280 n4145 n4146 n4144 VDD GND NOR2_X1
xU11281 n8430 n472 n4146 VDD GND NOR2_X1
xU11282 n8395 n287 n4145 VDD GND NOR2_X1
xU11283 \AES_Comp_ENCa/KrgX_65 n3063 n3056 VDD GND NOR2_X1
xU11284 n3064 n3065 n3063 VDD GND NOR2_X1
xU11285 n8428 n573 n3065 VDD GND NOR2_X1
xU11286 n8393 n233 n3064 VDD GND NOR2_X1
xU11287 n1579 n956 n1578 VDD GND NOR2_X1
xU11288 n1580 n1581 n1579 VDD GND NOR2_X1
xU11289 n8423 n143 n1581 VDD GND NOR2_X1
xU11290 n8389 n172 n1580 VDD GND NOR2_X1
xU11291 \AES_Comp_ENCa/KrgX_120 n1168 n1161 VDD GND NOR2_X1
xU11292 n1169 n1170 n1168 VDD GND NOR2_X1
xU11293 n8425 n659 n1170 VDD GND NOR2_X1
xU11294 n8391 n170 n1169 VDD GND NOR2_X1
xU11295 n5193 n842 n5192 VDD GND NOR2_X1
xU11296 n5194 n5195 n5193 VDD GND NOR2_X1
xU11297 n8432 n4965 n5195 VDD GND NOR2_X1
xU11298 n8397 n344 n5194 VDD GND NOR2_X1
xU11299 n1748 n951 n1747 VDD GND NOR2_X1
xU11300 n1749 n1750 n1748 VDD GND NOR2_X1
xU11301 n8424 n1751 n1750 VDD GND NOR2_X1
xU11302 n8391 n155 n1749 VDD GND NOR2_X1
xU11303 \AES_Comp_ENCa/KrgX_88 n2413 n2406 VDD GND NOR2_X1
xU11304 n2414 n2415 n2413 VDD GND NOR2_X1
xU11305 n8425 n547 n2415 VDD GND NOR2_X1
xU11306 n8391 n200 n2414 VDD GND NOR2_X1
xU11307 n1656 n953 n1655 VDD GND NOR2_X1
xU11308 n1657 n1658 n1656 VDD GND NOR2_X1
xU11309 n8424 n1073 n1658 VDD GND NOR2_X1
xU11310 n8389 n140 n1657 VDD GND NOR2_X1
xU11311 n4703 n884 n4702 VDD GND NOR2_X1
xU11312 n4704 n4705 n4703 VDD GND NOR2_X1
xU11313 n8430 n4706 n4705 VDD GND NOR2_X1
xU11314 n8396 n353 n4704 VDD GND NOR2_X1
xU11315 n1447 n961 n1446 VDD GND NOR2_X1
xU11316 n1448 n1449 n1447 VDD GND NOR2_X1
xU11317 n8424 n402 n1449 VDD GND NOR2_X1
xU11318 n8388 n145 n1448 VDD GND NOR2_X1
xU11319 \AES_Comp_ENCa/KrgX_40 n4048 n4041 VDD GND NOR2_X1
xU11320 n4049 n4050 n4048 VDD GND NOR2_X1
xU11321 n8430 n601 n4050 VDD GND NOR2_X1
xU11322 n8395 n258 n4049 VDD GND NOR2_X1
xU11323 n3986 n895 n3985 VDD GND NOR2_X1
xU11324 n3987 n3988 n3986 VDD GND NOR2_X1
xU11325 n8429 n606 n3988 VDD GND NOR2_X1
xU11326 n8395 n283 n3987 VDD GND NOR2_X1
xU11327 \AES_Comp_ENCa/KrgX_105 n1533 n1527 VDD GND NOR2_X1
xU11328 n1534 n1535 n1533 VDD GND NOR2_X1
xU11329 n8423 n399 n1535 VDD GND NOR2_X1
xU11330 n8389 n149 n1534 VDD GND NOR2_X1
xU11331 \AES_Comp_ENCa/KrgX_45 n3915 n3909 VDD GND NOR2_X1
xU11332 n3916 n3917 n3915 VDD GND NOR2_X1
xU11333 n8429 n603 n3917 VDD GND NOR2_X1
xU11334 n8395 n270 n3916 VDD GND NOR2_X1
xU11335 \AES_Comp_ENCa/KrgX_104 n1562 n1555 VDD GND NOR2_X1
xU11336 n1563 n1564 n1562 VDD GND NOR2_X1
xU11337 n8423 n396 n1564 VDD GND NOR2_X1
xU11338 n8389 n144 n1563 VDD GND NOR2_X1
xU11339 n3567 n912 n3566 VDD GND NOR2_X1
xU11340 n3568 n3569 n3567 VDD GND NOR2_X1
xU11341 n8428 n3570 n3569 VDD GND NOR2_X1
xU11342 n8394 n267 n3568 VDD GND NOR2_X1
xU11343 n2903 n921 n2902 VDD GND NOR2_X1
xU11344 n2904 n2905 n2903 VDD GND NOR2_X1
xU11345 n8427 n577 n2905 VDD GND NOR2_X1
xU11346 n8393 n229 n2904 VDD GND NOR2_X1
xU11347 \AES_Comp_ENCa/KrgX_96 n1872 n1865 VDD GND NOR2_X1
xU11348 n1873 n1874 n1872 VDD GND NOR2_X1
xU11349 n8425 n171 n1874 VDD GND NOR2_X1
xU11350 n8390 n138 n1873 VDD GND NOR2_X1
xU11351 \AES_Comp_ENCa/KrgX_32 n4351 n4345 VDD GND NOR2_X1
xU11352 n4352 n4353 n4351 VDD GND NOR2_X1
xU11353 n8430 n474 n4353 VDD GND NOR2_X1
xU11354 n8396 n256 n4352 VDD GND NOR2_X1
xU11355 n2996 n919 n2995 VDD GND NOR2_X1
xU11356 n2997 n2998 n2996 VDD GND NOR2_X1
xU11357 n8428 n576 n2998 VDD GND NOR2_X1
xU11358 n8393 n205 n2997 VDD GND NOR2_X1
xU11359 n2294 n945 n2293 VDD GND NOR2_X1
xU11360 n2295 n2296 n2294 VDD GND NOR2_X1
xU11361 n8424 n554 n2296 VDD GND NOR2_X1
xU11362 n8390 n232 n2295 VDD GND NOR2_X1
xU11363 \AES_Comp_ENCa/KrgX_49 n3821 n3814 VDD GND NOR2_X1
xU11364 n3822 n3823 n3821 VDD GND NOR2_X1
xU11365 n8429 n277 n3823 VDD GND NOR2_X1
xU11366 n8394 n263 n3822 VDD GND NOR2_X1
xU11367 n4999 n861 n4998 VDD GND NOR2_X1
xU11368 n5000 n5001 n4999 VDD GND NOR2_X1
xU11369 n8431 n4768 n5001 VDD GND NOR2_X1
xU11370 n8397 n345 n5000 VDD GND NOR2_X1
xU11371 \AES_Comp_ENCa/KrgX_112 n1364 n1357 VDD GND NOR2_X1
xU11372 n1365 n1366 n1364 VDD GND NOR2_X1
xU11373 n8423 n521 n1366 VDD GND NOR2_X1
xU11374 n8389 n169 n1365 VDD GND NOR2_X1
xU11375 \AES_Comp_ENCa/KrgX_81 n2582 n2575 VDD GND NOR2_X1
xU11376 n2583 n2584 n2582 VDD GND NOR2_X1
xU11377 n8426 n426 n2584 VDD GND NOR2_X1
xU11378 n8392 n220 n2583 VDD GND NOR2_X1
xU11379 n1280 n968 n1279 VDD GND NOR2_X1
xU11380 n1281 n1282 n1280 VDD GND NOR2_X1
xU11381 n8423 n1283 n1282 VDD GND NOR2_X1
xU11382 n8390 n177 n1281 VDD GND NOR2_X1
xU11383 n3760 n904 n3759 VDD GND NOR2_X1
xU11384 n3761 n3762 n3760 VDD GND NOR2_X1
xU11385 n8429 n3763 n3762 VDD GND NOR2_X1
xU11386 n8394 n291 n3761 VDD GND NOR2_X1
xU11387 \AES_Comp_ENCa/KrgX_16 n5077 n5070 VDD GND NOR2_X1
xU11388 n5078 n5079 n5077 VDD GND NOR2_X1
xU11389 n8431 n629 n5079 VDD GND NOR2_X1
xU11390 n8397 n341 n5078 VDD GND NOR2_X1
xU11391 \AES_Comp_ENCa/KrgX_117 n1237 n1231 VDD GND NOR2_X1
xU11392 n1238 n1239 n1237 VDD GND NOR2_X1
xU11393 n8425 n1240 n1239 VDD GND NOR2_X1
xU11394 n8389 n159 n1238 VDD GND NOR2_X1
xU11395 n3961 n896 n3960 VDD GND NOR2_X1
xU11396 n3962 n3963 n3961 VDD GND NOR2_X1
xU11397 n8429 n3728 n3963 VDD GND NOR2_X1
xU11398 n8395 n260 n3962 VDD GND NOR2_X1
xU11399 n1477 n960 n1476 VDD GND NOR2_X1
xU11400 n1478 n1479 n1477 VDD GND NOR2_X1
xU11401 n8423 n1480 n1479 VDD GND NOR2_X1
xU11402 n8388 n164 n1478 VDD GND NOR2_X1
xU11403 \AES_Comp_ENCa/KrgX_64 n3117 n3111 VDD GND NOR2_X1
xU11404 n3118 n3119 n3117 VDD GND NOR2_X1
xU11405 n8428 n2616 n3119 VDD GND NOR2_X1
xU11406 n8393 n198 n3118 VDD GND NOR2_X1
xU11407 \AES_Comp_ENCa/KrgX_97 n1817 n1810 VDD GND NOR2_X1
xU11408 n1818 n1819 n1817 VDD GND NOR2_X1
xU11409 n8424 n154 n1819 VDD GND NOR2_X1
xU11410 n8390 n139 n1818 VDD GND NOR2_X1
xU11411 \AES_Comp_ENCa/KrgX_0 n5587 n5581 VDD GND NOR2_X1
xU11412 n5588 n5589 n5587 VDD GND NOR2_X1
xU11413 n8426 n371 n5589 VDD GND NOR2_X1
xU11414 n8391 n313 n5588 VDD GND NOR2_X1
xU11415 Dout_E_89 n3019 n2865 VDD GND NAND2_X1
xU11416 n6632 n883 n6631 VDD GND NOR2_X1
xU11417 n6633 n8291 n6632 VDD GND NOR2_X1
xU11418 n6397 n8338 n6633 VDD GND AND2_X1
xU11419 n7116 n846 n7115 VDD GND NOR2_X1
xU11420 n7117 n8299 n7116 VDD GND NOR2_X1
xU11421 n6509 n8339 n7117 VDD GND AND2_X1
xU11422 n6696 n879 n6695 VDD GND NOR2_X1
xU11423 n6697 n8293 n6696 VDD GND NOR2_X1
xU11424 n6418 n8338 n6697 VDD GND AND2_X1
xU11425 n7228 n839 n7227 VDD GND NOR2_X1
xU11426 n7229 n8302 n7228 VDD GND NOR2_X1
xU11427 n6551 n8339 n7229 VDD GND AND2_X1
xU11428 n1892 n2069 n2038 VDD GND NAND2_X1
xU11429 n5599 n5676 n5669 VDD GND NAND2_X1
xU11430 n5563 n5741 n5737 VDD GND NAND2_X1
xU11431 n4386 n4439 n4431 VDD GND NAND2_X1
xU11432 n3147 n3208 n3197 VDD GND NAND2_X1
xU11433 n2149 n2199 n2191 VDD GND NAND2_X1
xU11434 n6794 n6844 n6835 VDD GND NAND2_X1
xU11435 n3129 n3272 n3256 VDD GND NAND2_X1
xU11436 n1881 n2119 n2112 VDD GND NAND2_X1
xU11437 n4362 n4605 n4598 VDD GND NAND2_X1
xU11438 n4625 n4671 n4661 VDD GND NAND2_X1
xU11439 n2141 n2188 n2176 VDD GND NAND2_X1
xU11440 n7012 n7091 n7063 VDD GND NAND2_X1
xU11441 n4459 n4511 n4499 VDD GND NAND2_X1
xU11442 n7242 n7315 n7291 VDD GND NAND2_X1
xU11443 n3392 n3446 n3426 VDD GND NAND2_X1
xU11444 n3155 n3204 n3180 VDD GND NAND2_X1
xU11445 \AES_Comp_ENCa/KrgX_5 n5343 n5337 VDD GND NOR2_X1
xU11446 n5344 n5345 n5343 VDD GND NOR2_X1
xU11447 n8432 n374 n5345 VDD GND NOR2_X1
xU11448 n8398 n339 n5344 VDD GND NOR2_X1
xU11449 \AES_Comp_ENCa/KrgX_6 n5320 n5313 VDD GND NOR2_X1
xU11450 n5321 n5322 n5320 VDD GND NOR2_X1
xU11451 n8432 n376 n5322 VDD GND NOR2_X1
xU11452 n8398 n315 n5321 VDD GND NOR2_X1
xU11453 n5781 n5833 n5809 VDD GND NAND2_X1
xU11454 Dout_E_46 n2000 n1968 VDD GND NAND2_X1
xU11455 n5782 n5846 n5826 VDD GND NAND2_X1
xU11456 n4393 n4424 n4418 VDD GND NAND2_X1
xU11457 n3316 n3354 n3340 VDD GND NAND2_X1
xU11458 n5546 n5904 n5896 VDD GND NAND2_X1
xU11459 n5618 n5685 n5668 VDD GND NAND2_X1
xU11460 n4474 n4506 n4497 VDD GND NAND2_X1
xU11461 n4361 n4607 n4593 VDD GND NAND2_X1
xU11462 n4539 n4667 n4658 VDD GND NAND2_X1
xU11463 n3385 n3440 n3423 VDD GND NAND2_X1
xU11464 n1884 n2122 n2108 VDD GND NAND2_X1
xU11465 n3148 n3212 n3188 VDD GND NAND2_X1
xU11466 n4359 n4587 n4582 VDD GND NAND2_X1
xU11467 n6795 n6841 n6832 VDD GND NAND2_X1
xU11468 n7464 n7513 n7503 VDD GND NAND2_X1
xU11469 n2156 n2185 n2177 VDD GND NAND2_X1
xU11470 n7020 n7089 n7059 VDD GND NAND2_X1
xU11471 \AES_Comp_ENCa/KrgX_30 n7531 n7494 VDD GND NAND2_X1
xU11472 n5897 n5871 n5890 VDD GND NAND2_X1
xU11473 n5613 n5597 n5544 VDD GND NAND2_X1
xU11474 n3242 n581 n2688 VDD GND NAND2_X1
xU11475 \AES_Comp_ENCa/KrgX_22 n6724 n6676 VDD GND NAND2_X1
xU11476 \AES_Comp_ENCa/KrgX_6 n7185 n7219 VDD GND NAND2_X1
xU11477 Dout_E_22 n4526 n4491 VDD GND NAND2_X1
xU11478 Dout_E_102 n3285 n3251 VDD GND NAND2_X1
xU11479 Dout_E_14 n3434 n3413 VDD GND NAND2_X1
xU11480 Dout_E_6 n2114 n2088 VDD GND NAND2_X1
xU11481 \AES_Comp_ENCa/KrgX_6 n7296 n7281 VDD GND NAND2_X1
xU11482 n1982 n1953 n1975 VDD GND NAND2_X1
xU11483 n588 n2918 n2917 VDD GND NOR2_X1
xU11484 n3309 n3362 n3334 VDD GND AND2_X1
xU11485 n6757 n6758 n6734 VDD GND NAND2_X1
xU11486 n1839 n1990 n1967 VDD GND AND2_X1
xU11487 n6995 n7065 n7047 VDD GND AND2_X1
xU11488 Dout_E_49 n3141 n3078 VDD GND NAND2_X1
xU11489 n3127 n3266 n3259 VDD GND NAND2_X1
xU11490 n5701 n5758 n5751 VDD GND NAND2_X1
xU11491 n7246 n7314 n7287 VDD GND NAND2_X1
xU11492 n3377 n3299 n3357 VDD GND NAND2_X1
xU11493 n3170 n3171 n2863 VDD GND AND2_X1
xU11494 n5929 n5493 n5914 VDD GND NAND2_X1
xU11495 Dout_E_38 n5671 n5665 VDD GND NAND2_X1
xU11496 Dout_E_118 n5919 n5912 VDD GND NAND2_X1
xU11497 \AES_Comp_ENCa/KrgX_1 n7236 n7206 VDD GND NAND2_X1
xU11498 Dout_E_110 n4442 n4412 VDD GND NAND2_X1
xU11499 Dout_E_54 n3198 n3186 VDD GND NAND2_X1
xU11500 Dout_E_86 n2202 n2172 VDD GND NAND2_X1
xU11501 \AES_Comp_ENCa/KrgX_30 n7410 n7378 VDD GND NAND2_X1
xU11502 n4617 n4367 n4583 VDD GND NAND2_X1
xU11503 n5767 n5487 n5752 VDD GND NAND2_X1
xU11504 Dout_E_94 n3349 n3344 VDD GND NAND2_X1
xU11505 Dout_E_94 n3047 n2720 VDD GND NAND2_X1
xU11506 Dout_E_78 n5755 n5749 VDD GND NAND2_X1
xU11507 Dout_E_78 n5503 n5432 VDD GND NAND2_X1
xU11508 n4549 n482 n4325 VDD GND NAND2_X1
xU11509 Dout_E_30 n5827 n5819 VDD GND NAND2_X1
xU11510 n6961 n6962 n6928 VDD GND NAND2_X1
xU11511 n5682 n5683 n5673 VDD GND NAND2_X1
xU11512 n5616 n388 n5683 VDD GND OR2_X1
xU11513 n5616 n391 n5682 VDD GND NAND2_X1
xU11514 n6864 n6865 n6834 VDD GND NAND2_X1
xU11515 n6753 n857 n6865 VDD GND OR2_X1
xU11516 n6753 n863 n6864 VDD GND NAND2_X1
xU11517 n4531 n4532 n4500 VDD GND NAND2_X1
xU11518 n4334 n303 n4532 VDD GND OR2_X1
xU11519 n4334 n4515 n4531 VDD GND NAND2_X1
xU11520 Dout_E_70 n4601 n4595 VDD GND NAND2_X1
xU11521 n7409 n7410 n7377 VDD GND NAND2_X1
xU11522 n4251 n4252 n4157 VDD GND NAND2_X1
xU11523 n3007 n3008 n2916 VDD GND NAND2_X1
xU11524 n4264 n4265 n4183 VDD GND NAND2_X1
xU11525 n1761 n1762 n1668 VDD GND NAND2_X1
xU11526 n4283 n4284 n4173 VDD GND NAND2_X1
xU11527 n7184 n7185 n7148 VDD GND NAND2_X1
xU11528 n3029 n3030 n2950 VDD GND NAND2_X1
xU11529 n5474 n5475 n5380 VDD GND NAND2_X1
xU11530 n1782 n1783 n1712 VDD GND NAND2_X1
xU11531 n5502 n5503 n5425 VDD GND NAND2_X1
xU11532 n6723 n6724 n6684 VDD GND NAND2_X1
xU11533 Dout_E_126 n2071 n2053 VDD GND NAND2_X1
xU11534 n1773 n1774 n1683 VDD GND NAND2_X1
xU11535 n3038 n3039 n2932 VDD GND NAND2_X1
xU11536 n4291 n4292 n4201 VDD GND NAND2_X1
xU11537 n1794 n1795 n1693 VDD GND NAND2_X1
xU11538 Dout_E_113 n5853 n5548 VDD GND AND2_X1
xU11539 Dout_E_41 n1935 n1843 VDD GND AND2_X1
xU11540 Dout_E_17 n4456 n4328 VDD GND AND2_X1
xU11541 n4432 n4320 n4413 VDD GND AND2_X1
xU11542 \AES_Comp_ENCa/KrgX_17 n6790 n6755 VDD GND AND2_X1
xU11543 Dout_E_33 n5609 n5596 VDD GND AND2_X1
xU11544 n3022 n3370 n3345 VDD GND AND2_X1
xU11545 n4382 n4450 n4419 VDD GND AND2_X1
xU11546 n4541 n4612 n4596 VDD GND AND2_X1
xU11547 n4273 n4689 n4659 VDD GND AND2_X1
xU11548 n2145 n2206 n2178 VDD GND AND2_X1
xU11549 n1804 n2063 n2050 VDD GND AND2_X1
xU11550 n1911 n2130 n2109 VDD GND AND2_X1
xU11551 n1857 n2054 n2039 VDD GND AND2_X1
xU11552 n5856 n5902 n5891 VDD GND AND2_X1
xU11553 n1938 n1986 n1974 VDD GND AND2_X1
xU11554 n7462 n7535 n7504 VDD GND AND2_X1
xU11555 n5598 n5658 n5650 VDD GND AND2_X1
xU11556 Dout_E_81 n2137 n1831 VDD GND AND2_X1
xU11557 Dout_E_57 n4270 n4106 VDD GND AND2_X1
xU11558 Dout_E_9 n3380 n3093 VDD GND AND2_X1
xU11559 Dout_E_121 n1801 n1615 VDD GND AND2_X1
xU11560 n6793 n6866 n6833 VDD GND AND2_X1
xU11561 n4309 n4599 n4594 VDD GND AND2_X1
xU11562 \AES_Comp_ENCa/KrgX_14 n6962 n6999 VDD GND AND2_X1
xU11563 n2192 n1830 n2173 VDD GND AND2_X1
xU11564 n3372 n3373 n3348 VDD GND NAND2_X1
xU11565 n562 n3375 n3372 VDD GND NAND2_X1
xU11566 n3374 Dout_E_89 n3373 VDD GND NAND2_X1
xU11567 n5925 n5926 n5918 VDD GND NAND2_X1
xU11568 n5927 Dout_E_113 n5926 VDD GND NAND2_X1
xU11569 n645 n652 n5925 VDD GND NAND2_X1
xU11570 Dout_E_54 n3039 n2940 VDD GND AND2_X1
xU11571 Dout_E_110 n4265 n4191 VDD GND AND2_X1
xU11572 Dout_E_86 n1783 n1719 VDD GND AND2_X1
xU11573 Dout_E_118 n5511 n5408 VDD GND AND2_X1
xU11574 Dout_E_38 n5475 n5388 VDD GND AND2_X1
xU11575 Dout_E_46 n1795 n1701 VDD GND AND2_X1
xU11576 n358 n5800 n5786 VDD GND NAND2_X1
xU11577 Dout_E_62 n4284 n3952 VDD GND AND2_X1
xU11578 n5491 n5844 n5820 VDD GND AND2_X1
xU11579 n7216 n7305 n7295 VDD GND AND2_X1
xU11580 n5860 n5923 n5913 VDD GND AND2_X1
xU11581 n3162 n3217 n3189 VDD GND AND2_X1
xU11582 n4533 n4463 n4498 VDD GND AND2_X1
xU11583 n3458 n3399 n3424 VDD GND AND2_X1
xU11584 n3293 n3137 n3260 VDD GND AND2_X1
xU11585 n2008 n1942 n1976 VDD GND AND2_X1
xU11586 n5762 n5697 n5750 VDD GND AND2_X1
xU11587 n7087 n7016 n7082 VDD GND AND2_X1
xU11588 n7288 n7245 n7280 VDD GND AND2_X1
xU11589 n6971 n7083 n7060 VDD GND AND2_X1
xU11590 n3134 n3295 n3265 VDD GND AND2_X1
xU11591 Dout_E_30 n5519 n5184 VDD GND AND2_X1
xU11592 n5775 n5838 n5810 VDD GND AND2_X1
xU11593 n7463 n7517 n7506 VDD GND AND2_X1
xU11594 n4378 n4428 n4417 VDD GND AND2_X1
xU11595 n7238 n7307 n7282 VDD GND AND2_X1
xU11596 n1897 n2057 n2033 VDD GND AND2_X1
xU11597 n5536 n5661 n5655 VDD GND AND2_X1
xU11598 n3018 n3460 n3439 VDD GND AND2_X1
xU11599 Dout_E_126 n1774 n1469 VDD GND AND2_X1
xU11600 Dout_E_70 n4252 n4165 VDD GND AND2_X1
xU11601 Dout_E_6 n1762 n1675 VDD GND AND2_X1
xU11602 Dout_E_102 n3008 n2923 VDD GND AND2_X1
xU11603 n5680 n5629 n5666 VDD GND AND2_X1
xU11604 n4694 n4695 n4660 VDD GND NAND2_X1
xU11605 n4628 n460 n4695 VDD GND OR2_X1
xU11606 n4628 n464 n4694 VDD GND NAND2_X1
xU11607 n2212 n2213 n2175 VDD GND NAND2_X1
xU11608 n1838 n539 n2213 VDD GND OR2_X1
xU11609 n1838 n2193 n2212 VDD GND NAND2_X1
xU11610 n2128 n2129 n2111 VDD GND NAND2_X1
xU11611 n1924 n190 n2129 VDD GND OR2_X1
xU11612 n1924 n193 n2128 VDD GND NAND2_X1
xU11613 n4614 n4615 n4600 VDD GND NAND2_X1
xU11614 n4553 n485 n4615 VDD GND OR2_X1
xU11615 n4553 n491 n4614 VDD GND NAND2_X1
xU11616 n7292 n7293 n7275 VDD GND NAND2_X1
xU11617 n7210 n825 n7293 VDD GND OR2_X1
xU11618 n7210 n828 n7292 VDD GND NAND2_X1
xU11619 n7092 n7093 n7080 VDD GND NAND2_X1
xU11620 n6988 n840 n7093 VDD GND OR2_X1
xU11621 n6988 n843 n7092 VDD GND NAND2_X1
xU11622 n3291 n3292 n3255 VDD GND NAND2_X1
xU11623 n3224 n593 n3292 VDD GND OR2_X1
xU11624 n3224 n596 n3291 VDD GND NAND2_X1
xU11625 n5764 n5765 n5754 VDD GND NAND2_X1
xU11626 n5572 n513 n5765 VDD GND OR2_X1
xU11627 n5572 n5742 n5764 VDD GND NAND2_X1
xU11628 n4448 n4449 n4416 VDD GND NAND2_X1
xU11629 n4319 n618 n4449 VDD GND OR2_X1
xU11630 n4319 n624 n4448 VDD GND NAND2_X1
xU11631 n3222 n3223 n3179 VDD GND NAND2_X1
xU11632 n3084 n434 n3223 VDD GND OR2_X1
xU11633 n3084 n439 n3222 VDD GND NAND2_X1
xU11634 n3456 n3457 n3425 VDD GND NAND2_X1
xU11635 n3099 n245 n3457 VDD GND OR2_X1
xU11636 n3099 n251 n3456 VDD GND NAND2_X1
xU11637 n2073 n2074 n2056 VDD GND NAND2_X1
xU11638 n1901 n669 n2074 VDD GND OR2_X1
xU11639 n1901 n676 n2073 VDD GND NAND2_X1
xU11640 n5656 n5601 n5649 VDD GND AND2_X1
xU11641 Dout_E_22 n4292 n4209 VDD GND AND2_X1
xU11642 Dout_E_14 n3030 n2958 VDD GND AND2_X1
xU11643 n7537 n7419 n7512 VDD GND AND2_X1
xU11644 n4452 n4277 n4423 VDD GND AND2_X1
xU11645 n4691 n4368 n4666 VDD GND AND2_X1
xU11646 n6868 n6737 n6840 VDD GND AND2_X1
xU11647 n3219 n3024 n3211 VDD GND AND2_X1
xU11648 n2208 n1787 n2184 VDD GND AND2_X1
xU11649 n2065 n2012 n2037 VDD GND AND2_X1
xU11650 n2132 n2075 n2121 VDD GND AND2_X1
xU11651 n7311 n7190 n7279 VDD GND AND2_X1
xU11652 n4535 n4279 n4505 VDD GND AND2_X1
xU11653 n2010 n1800 n1981 VDD GND AND2_X1
xU11654 n6992 n6993 n6973 VDD GND AND2_X1
xU11655 n7213 n7214 n7192 VDD GND AND2_X1
xU11656 n7440 n871 n7421 VDD GND AND2_X1
xU11657 n5788 n5780 n5327 VDD GND AND2_X1
xU11658 n8253 n8254 n1973 VDD GND NOR2_X1
xU11659 n1841 n414 n8253 VDD GND AND2_X1
xU11660 n1841 n411 n8254 VDD GND NOR2_X1
xU11661 n4175 n4176 n4174 VDD GND NAND2_X1
xU11662 n6686 n6687 n6685 VDD GND NAND2_X1
xU11663 n2934 n430 n2933 VDD GND NOR2_X1
xU11664 n2935 n430 VDD GND INV_X1
xU11665 n4854 n4855 n7948 VDD GND NAND2_X1
xU11666 n4876 n4877 n4854 VDD GND NOR2_X1
xU11667 n4856 n4857 n4855 VDD GND NOR2_X1
xU11668 n8368 n362 n4877 VDD GND NOR2_X1
xU11669 n5157 n5158 n7961 VDD GND NAND2_X1
xU11670 n5186 n5187 n5157 VDD GND NOR2_X1
xU11671 n5159 n5160 n5158 VDD GND NOR2_X1
xU11672 n8369 n252 n5187 VDD GND NOR2_X1
xU11673 n5456 n5457 n7971 VDD GND NAND2_X1
xU11674 n5521 n5522 n5456 VDD GND NOR2_X1
xU11675 n5458 n5459 n5457 VDD GND NOR2_X1
xU11676 n191 n8357 n5522 VDD GND NOR2_X1
xU11677 n1398 n1399 n7863 VDD GND NAND2_X1
xU11678 n1418 n1419 n1398 VDD GND NOR2_X1
xU11679 n1400 n1401 n1399 VDD GND NOR2_X1
xU11680 n8361 n627 n1419 VDD GND NOR2_X1
xU11681 n2823 n2824 n7902 VDD GND NAND2_X1
xU11682 n2842 n2843 n2823 VDD GND NOR2_X1
xU11683 n2825 n2826 n2824 VDD GND NOR2_X1
xU11684 n8364 n495 n2843 VDD GND NOR2_X1
xU11685 n1179 n1180 n7854 VDD GND NAND2_X1
xU11686 n1202 n1203 n1179 VDD GND NOR2_X1
xU11687 n1181 n1182 n1180 VDD GND NOR2_X1
xU11688 n8360 n656 n1203 VDD GND NOR2_X1
xU11689 n1250 n1251 n7857 VDD GND NAND2_X1
xU11690 n1273 n1274 n1250 VDD GND NOR2_X1
xU11691 n1252 n1253 n1251 VDD GND NOR2_X1
xU11692 n8361 n653 n1274 VDD GND NOR2_X1
xU11693 n2696 n2697 n7897 VDD GND NAND2_X1
xU11694 n2724 n2725 n2696 VDD GND NOR2_X1
xU11695 n2698 n2699 n2697 VDD GND NOR2_X1
xU11696 n8364 n517 n2725 VDD GND NOR2_X1
xU11697 n3781 n3782 n7923 VDD GND NAND2_X1
xU11698 n3809 n3810 n3781 VDD GND NOR2_X1
xU11699 n3783 n3784 n3782 VDD GND NOR2_X1
xU11700 n8366 n436 n3810 VDD GND NOR2_X1
xU11701 n1597 n1598 n7871 VDD GND NAND2_X1
xU11702 n1619 n1620 n1597 VDD GND NOR2_X1
xU11703 n1599 n1600 n1598 VDD GND NOR2_X1
xU11704 n8362 n599 n1620 VDD GND NOR2_X1
xU11705 n2475 n2476 n7888 VDD GND NAND2_X1
xU11706 n2496 n2497 n2475 VDD GND NOR2_X1
xU11707 n2477 n2478 n2476 VDD GND NOR2_X1
xU11708 n544 n8360 n2497 VDD GND NOR2_X1
xU11709 n7574 n7575 n7573 VDD GND NAND2_X1
xU11710 n133 n981 n7575 VDD GND NAND2_X1
xU11711 BSY_E n813 n7574 VDD GND NAND2_X1
xU11712 RSTn n8330 n7570 VDD GND NAND2_X1
xU11713 n6767 n6768 n6656 VDD GND NAND2_X1
xU11714 \AES_Comp_ENCa/Rrg_8 \AES_Comp_ENCa/Rrg_7 n6768 VDD GND NOR2_X1
xU11715 n6625 n817 n6767 VDD GND NOR2_X1
xU11716 n6787 n811 n6625 VDD GND NAND2_X1
xU11717 \AES_Comp_ENCa/Rrg_6 \AES_Comp_ENCa/Rrg_5 n6787 VDD GND NOR2_X1
xU11718 n6786 \AES_Comp_ENCa/Rrg_8 n6680 VDD GND NAND2_X1
xU11719 \AES_Comp_ENCa/Rrg_7 n6625 n6786 VDD GND NOR2_X1
xU11720 n6789 n813 n6704 VDD GND NAND2_X1
xU11721 \AES_Comp_ENCa/Rrg_2 \AES_Comp_ENCa/Rrg_1 n6789 VDD GND NOR2_X1
xU11722 n6704 n814 n6703 VDD GND NOR2_X1
xU11723 \AES_Comp_ENCa/Rrg_5 n6641 n6640 VDD GND NOR2_X1
xU11724 n7567 RSTn n8112 VDD GND NAND2_X1
xU11725 n7568 n7569 n7567 VDD GND NOR2_X1
xU11726 n813 n7570 n7569 VDD GND NOR2_X1
xU11727 \AES_Comp_ENCa/Rrg_9 n7546 n7568 VDD GND AND2_X1
xU11728 n6625 n816 n6624 VDD GND NOR2_X1
xU11729 n6788 n812 n6641 VDD GND NAND2_X1
xU11730 \AES_Comp_ENCa/Rrg_4 \AES_Comp_ENCa/Rrg_3 n6788 VDD GND NOR2_X1
xU11731 n812 n814 n6681 VDD GND NAND2_X1
xU11732 n7452 n981 n5931 VDD GND NOR2_X1
xU11733 BSY_E n7452 n5935 VDD GND NOR2_X1
xU11734 n753 n8418 n6326 VDD GND NOR2_X1
xU11735 n745 n8417 n6382 VDD GND NOR2_X1
xU11736 n713 n8415 n6606 VDD GND NOR2_X1
xU11737 n749 n8418 n6354 VDD GND NOR2_X1
xU11738 n786 n8418 n6095 VDD GND NOR2_X1
xU11739 n754 n8418 n6319 VDD GND NOR2_X1
xU11740 n746 n8418 n6375 VDD GND NOR2_X1
xU11741 n755 n8418 n6312 VDD GND NOR2_X1
xU11742 n748 n8418 n6361 VDD GND NOR2_X1
xU11743 n750 n8418 n6347 VDD GND NOR2_X1
xU11744 n747 n8418 n6368 VDD GND NOR2_X1
xU11745 n751 n8418 n6340 VDD GND NOR2_X1
xU11746 n752 n8418 n6333 VDD GND NOR2_X1
xU11747 n720 n8415 n6557 VDD GND NOR2_X1
xU11748 n742 n8417 n6403 VDD GND NOR2_X1
xU11749 n736 n8417 n6445 VDD GND NOR2_X1
xU11750 n733 n8416 n6466 VDD GND NOR2_X1
xU11751 n725 n8416 n6522 VDD GND NOR2_X1
xU11752 n719 n8415 n6564 VDD GND NOR2_X1
xU11753 n743 n8417 n6396 VDD GND NOR2_X1
xU11754 n734 n8417 n6459 VDD GND NOR2_X1
xU11755 n728 n8416 n6501 VDD GND NOR2_X1
xU11756 n715 n8415 n6592 VDD GND NOR2_X1
xU11757 n739 n8417 n6424 VDD GND NOR2_X1
xU11758 n735 n8417 n6452 VDD GND NOR2_X1
xU11759 n727 n8416 n6508 VDD GND NOR2_X1
xU11760 n718 n8415 n6571 VDD GND NOR2_X1
xU11761 n744 n8417 n6389 VDD GND NOR2_X1
xU11762 n731 n8416 n6480 VDD GND NOR2_X1
xU11763 n724 n8416 n6529 VDD GND NOR2_X1
xU11764 n726 n8416 n6515 VDD GND NOR2_X1
xU11765 n716 n8415 n6585 VDD GND NOR2_X1
xU11766 n741 n8417 n6410 VDD GND NOR2_X1
xU11767 n740 n8417 n6417 VDD GND NOR2_X1
xU11768 n732 n8416 n6473 VDD GND NOR2_X1
xU11769 n723 n8416 n6536 VDD GND NOR2_X1
xU11770 n714 n8415 n6599 VDD GND NOR2_X1
xU11771 n738 n8417 n6431 VDD GND NOR2_X1
xU11772 n730 n8416 n6487 VDD GND NOR2_X1
xU11773 n722 n8416 n6543 VDD GND NOR2_X1
xU11774 n717 n8415 n6578 VDD GND NOR2_X1
xU11775 n737 n8417 n6438 VDD GND NOR2_X1
xU11776 n729 n8416 n6494 VDD GND NOR2_X1
xU11777 n721 n8415 n6550 VDD GND NOR2_X1
xU11778 n3685 n8345 n3683 VDD GND NOR2_X1
xU11779 n3906 n8344 n3904 VDD GND NOR2_X1
xU11780 n4922 n8342 n4920 VDD GND NOR2_X1
xU11781 n3710 n8345 n3708 VDD GND NOR2_X1
xU11782 n3883 n8344 n3881 VDD GND NOR2_X1
xU11783 n3662 n8345 n3660 VDD GND NOR2_X1
xU11784 n3640 n8345 n3638 VDD GND NOR2_X1
xU11785 n3731 n8345 n3729 VDD GND NOR2_X1
xU11786 n4945 n8342 n4943 VDD GND NOR2_X1
xU11787 n4774 n8343 n4772 VDD GND NOR2_X1
xU11788 n4109 n8344 n4107 VDD GND NOR2_X1
xU11789 n3755 n8345 n3753 VDD GND NOR2_X1
xU11790 n4994 n8342 n4992 VDD GND NOR2_X1
xU11791 n5363 n8341 n5361 VDD GND NOR2_X1
xU11792 n4753 n8343 n4751 VDD GND NOR2_X1
xU11793 n4082 n8344 n4080 VDD GND NOR2_X1
xU11794 n5235 n8341 n5233 VDD GND NOR2_X1
xU11795 n3956 n8344 n3954 VDD GND NOR2_X1
xU11796 n5112 n8342 n5110 VDD GND NOR2_X1
xU11797 n5334 n8341 n5332 VDD GND NOR2_X1
xU11798 n3811 n8345 n3809 VDD GND NOR2_X1
xU11799 n4968 n8342 n4966 VDD GND NOR2_X1
xU11800 n5188 n8342 n5186 VDD GND NOR2_X1
xU11801 n5136 n8342 n5134 VDD GND NOR2_X1
xU11802 n5288 n8341 n5286 VDD GND NOR2_X1
xU11803 n5156 n8342 n5154 VDD GND NOR2_X1
xU11804 n5265 n8341 n5263 VDD GND NOR2_X1
xU11805 n5436 n8341 n5434 VDD GND NOR2_X1
xU11806 n4853 n8343 n4851 VDD GND NOR2_X1
xU11807 n4799 n8343 n4797 VDD GND NOR2_X1
xU11808 n4825 n8343 n4823 VDD GND NOR2_X1
xU11809 n4898 n8343 n4896 VDD GND NOR2_X1
xU11810 n4139 n8344 n4137 VDD GND NOR2_X1
xU11811 n5041 n8342 n5039 VDD GND NOR2_X1
xU11812 n4212 n8344 n4210 VDD GND NOR2_X1
xU11813 n5210 n8341 n5208 VDD GND NOR2_X1
xU11814 n5523 n8341 n5521 VDD GND NOR2_X1
xU11815 n4297 n8343 n4295 VDD GND NOR2_X1
xU11816 n5578 n8341 n5576 VDD GND NOR2_X1
xU11817 n4878 n8343 n4876 VDD GND NOR2_X1
xU11818 n4728 n8343 n4726 VDD GND NOR2_X1
xU11819 n4342 n8343 n4340 VDD GND NOR2_X1
xU11820 n4059 n8344 n4057 VDD GND NOR2_X1
xU11821 n4007 n8344 n4005 VDD GND NOR2_X1
xU11822 n3617 n8345 n3615 VDD GND NOR2_X1
xU11823 n3926 n8344 n3924 VDD GND NOR2_X1
xU11824 n4038 n8344 n4036 VDD GND NOR2_X1
xU11825 n3589 n8345 n3587 VDD GND NOR2_X1
xU11826 n5310 n8341 n5308 VDD GND NOR2_X1
xU11827 n4698 n8343 n4696 VDD GND NOR2_X1
xU11828 n3839 n8345 n3837 VDD GND NOR2_X1
xU11829 n5017 n8342 n5015 VDD GND NOR2_X1
xU11830 n3859 n8345 n3857 VDD GND NOR2_X1
xU11831 n5067 n8342 n5065 VDD GND NOR2_X1
xU11832 n3780 n8345 n3778 VDD GND NOR2_X1
xU11833 n5089 n8342 n5087 VDD GND NOR2_X1
xU11834 n3981 n8344 n3979 VDD GND NOR2_X1
xU11835 n5455 n8341 n5453 VDD GND NOR2_X1
xU11836 n4233 n8343 n4231 VDD GND NOR2_X1
xU11837 n5934 n8341 n5932 VDD GND NOR2_X1
xU11838 n682 n8418 n7443 VDD GND NOR2_X1
xU11839 n688 n8413 n7330 VDD GND NOR2_X1
xU11840 n710 n8415 n6661 VDD GND NOR2_X1
xU11841 n704 n8414 n6886 VDD GND NOR2_X1
xU11842 n701 n8414 n6932 VDD GND NOR2_X1
xU11843 n693 n8413 n7152 VDD GND NOR2_X1
xU11844 n687 n8413 n7342 VDD GND NOR2_X1
xU11845 n711 n8415 n6642 VDD GND NOR2_X1
xU11846 n702 n8414 n6911 VDD GND NOR2_X1
xU11847 n696 n8413 n7110 VDD GND NOR2_X1
xU11848 n707 n8414 n6738 VDD GND NOR2_X1
xU11849 n703 n8414 n6898 VDD GND NOR2_X1
xU11850 n695 n8413 n7122 VDD GND NOR2_X1
xU11851 n686 n8413 n7357 VDD GND NOR2_X1
xU11852 n712 n8415 n6626 VDD GND NOR2_X1
xU11853 n699 n8414 n6974 VDD GND NOR2_X1
xU11854 n692 n8413 n7163 VDD GND NOR2_X1
xU11855 n694 n8413 n7133 VDD GND NOR2_X1
xU11856 n709 n8414 n6690 VDD GND NOR2_X1
xU11857 n708 n8414 n6706 VDD GND NOR2_X1
xU11858 n700 n8414 n6944 VDD GND NOR2_X1
xU11859 n691 n8413 n7193 VDD GND NOR2_X1
xU11860 n706 n8414 n6769 VDD GND NOR2_X1
xU11861 n698 n8414 n7001 VDD GND NOR2_X1
xU11862 n690 n8413 n7222 VDD GND NOR2_X1
xU11863 n705 n8414 n6870 VDD GND NOR2_X1
xU11864 n697 n8413 n7094 VDD GND NOR2_X1
xU11865 n689 n8413 n7316 VDD GND NOR2_X1
xU11866 n681 n8402 n7542 VDD GND NOR2_X1
xU11867 n7544 n7545 n8102 VDD GND NAND2_X1
xU11868 n131 \AES_Comp_ENCa/Rrg_9 n7544 VDD GND NAND2_X1
xU11869 n7546 \AES_Comp_ENCa/Rrg_8 n7545 VDD GND NAND2_X1
xU11870 n7547 n7548 n8103 VDD GND NAND2_X1
xU11871 n131 \AES_Comp_ENCa/Rrg_8 n7547 VDD GND NAND2_X1
xU11872 n7546 \AES_Comp_ENCa/Rrg_7 n7548 VDD GND NAND2_X1
xU11873 n7549 n7550 n8104 VDD GND NAND2_X1
xU11874 n131 \AES_Comp_ENCa/Rrg_7 n7549 VDD GND NAND2_X1
xU11875 n7546 \AES_Comp_ENCa/Rrg_6 n7550 VDD GND NAND2_X1
xU11876 n7551 n7552 n8105 VDD GND NAND2_X1
xU11877 n131 \AES_Comp_ENCa/Rrg_6 n7551 VDD GND NAND2_X1
xU11878 n7546 \AES_Comp_ENCa/Rrg_5 n7552 VDD GND NAND2_X1
xU11879 n7553 n7554 n8106 VDD GND NAND2_X1
xU11880 n131 \AES_Comp_ENCa/Rrg_5 n7553 VDD GND NAND2_X1
xU11881 n7546 \AES_Comp_ENCa/Rrg_4 n7554 VDD GND NAND2_X1
xU11882 n7555 n7556 n8107 VDD GND NAND2_X1
xU11883 n131 \AES_Comp_ENCa/Rrg_4 n7555 VDD GND NAND2_X1
xU11884 n7546 \AES_Comp_ENCa/Rrg_3 n7556 VDD GND NAND2_X1
xU11885 n7557 n7558 n8108 VDD GND NAND2_X1
xU11886 n131 \AES_Comp_ENCa/Rrg_3 n7557 VDD GND NAND2_X1
xU11887 n7546 \AES_Comp_ENCa/Rrg_2 n7558 VDD GND NAND2_X1
xU11888 n7571 n7572 n8113 VDD GND NAND2_X1
xU11889 n131 \AES_Comp_ENCa/Rrg_2 n7571 VDD GND NAND2_X1
xU11890 n7546 \AES_Comp_ENCa/Rrg_1 n7572 VDD GND NAND2_X1
xU11891 n7559 n7560 n8109 VDD GND NAND2_X1
xU11892 n131 \AES_Comp_ENCa/Rrg_1 n7559 VDD GND NAND2_X1
xU11893 n7546 \AES_Comp_ENCa/Rrg_0 n7560 VDD GND NAND2_X1
xU11894 n5931 \AES_Comp_ENCa/Rrg_0 n989 VDD GND NAND2_X1
xU11895 n5931 n813 n991 VDD GND NAND2_X1
xU11896 n1053 n8351 n1051 VDD GND NOR2_X1
xU11897 n1081 n8351 n1079 VDD GND NOR2_X1
xU11898 n1106 n8351 n1104 VDD GND NOR2_X1
xU11899 n1158 n8351 n1156 VDD GND NOR2_X1
xU11900 n1032 n8351 n1030 VDD GND NOR2_X1
xU11901 n1134 n8351 n1132 VDD GND NOR2_X1
xU11902 n1178 n8351 n1176 VDD GND NOR2_X1
xU11903 n1008 n8351 n1005 VDD GND NOR2_X1
xU11904 n957 n8286 n6105 VDD GND NOR2_X1
xU11905 n925 n8289 n6329 VDD GND NOR2_X1
xU11906 n965 n8286 n6049 VDD GND NOR2_X1
xU11907 n933 n8288 n6273 VDD GND NOR2_X1
xU11908 n973 n8286 n5993 VDD GND NOR2_X1
xU11909 n941 n8288 n6217 VDD GND NOR2_X1
xU11910 n949 n8287 n6161 VDD GND NOR2_X1
xU11911 n917 n8287 n6385 VDD GND NOR2_X1
xU11912 n953 n8287 n6133 VDD GND NOR2_X1
xU11913 n921 n8289 n6357 VDD GND NOR2_X1
xU11914 n958 n8286 n6098 VDD GND NOR2_X1
xU11915 n926 n8289 n6322 VDD GND NOR2_X1
xU11916 n966 n8286 n6042 VDD GND NOR2_X1
xU11917 n934 n8288 n6266 VDD GND NOR2_X1
xU11918 n974 n8290 n5986 VDD GND NOR2_X1
xU11919 n942 n8288 n6210 VDD GND NOR2_X1
xU11920 n950 n8287 n6154 VDD GND NOR2_X1
xU11921 n918 n8286 n6378 VDD GND NOR2_X1
xU11922 n959 n8286 n6091 VDD GND NOR2_X1
xU11923 n927 n8289 n6315 VDD GND NOR2_X1
xU11924 n968 n8286 n6028 VDD GND NOR2_X1
xU11925 n936 n8288 n6252 VDD GND NOR2_X1
xU11926 n977 n8289 n5965 VDD GND NOR2_X1
xU11927 n945 n8287 n6189 VDD GND NOR2_X1
xU11928 n952 n8287 n6140 VDD GND NOR2_X1
xU11929 n920 n8288 n6364 VDD GND NOR2_X1
xU11930 n960 n8286 n6084 VDD GND NOR2_X1
xU11931 n928 n8289 n6308 VDD GND NOR2_X1
xU11932 n967 n8286 n6035 VDD GND NOR2_X1
xU11933 n935 n8288 n6259 VDD GND NOR2_X1
xU11934 n980 n8288 n5943 VDD GND NOR2_X1
xU11935 n948 n8287 n6168 VDD GND NOR2_X1
xU11936 n954 n8287 n6126 VDD GND NOR2_X1
xU11937 n922 n8289 n6350 VDD GND NOR2_X1
xU11938 n963 n8286 n6063 VDD GND NOR2_X1
xU11939 n931 n8289 n6287 VDD GND NOR2_X1
xU11940 n971 n8287 n6007 VDD GND NOR2_X1
xU11941 n939 n8288 n6231 VDD GND NOR2_X1
xU11942 n975 n8286 n5979 VDD GND NOR2_X1
xU11943 n943 n8288 n6203 VDD GND NOR2_X1
xU11944 n951 n8287 n6147 VDD GND NOR2_X1
xU11945 n919 n8289 n6371 VDD GND NOR2_X1
xU11946 n964 n8286 n6056 VDD GND NOR2_X1
xU11947 n932 n8289 n6280 VDD GND NOR2_X1
xU11948 n970 n8290 n6014 VDD GND NOR2_X1
xU11949 n938 n8288 n6238 VDD GND NOR2_X1
xU11950 n979 n8289 n5951 VDD GND NOR2_X1
xU11951 n947 n8287 n6175 VDD GND NOR2_X1
xU11952 n955 n8287 n6119 VDD GND NOR2_X1
xU11953 n923 n8289 n6343 VDD GND NOR2_X1
xU11954 n961 n8286 n6077 VDD GND NOR2_X1
xU11955 n929 n8289 n6301 VDD GND NOR2_X1
xU11956 n972 n8288 n6000 VDD GND NOR2_X1
xU11957 n940 n8288 n6224 VDD GND NOR2_X1
xU11958 n978 n8287 n5958 VDD GND NOR2_X1
xU11959 n946 n8287 n6182 VDD GND NOR2_X1
xU11960 n956 n8287 n6112 VDD GND NOR2_X1
xU11961 n924 n8289 n6336 VDD GND NOR2_X1
xU11962 n914 n8288 n6406 VDD GND NOR2_X1
xU11963 n969 n8286 n6021 VDD GND NOR2_X1
xU11964 n937 n8288 n6245 VDD GND NOR2_X1
xU11965 n915 n8290 n6399 VDD GND NOR2_X1
xU11966 n911 n8290 n6427 VDD GND NOR2_X1
xU11967 n916 n8287 n6392 VDD GND NOR2_X1
xU11968 n962 n8286 n6070 VDD GND NOR2_X1
xU11969 n930 n8289 n6294 VDD GND NOR2_X1
xU11970 n913 n8286 n6413 VDD GND NOR2_X1
xU11971 n976 n8290 n5972 VDD GND NOR2_X1
xU11972 n944 n8288 n6196 VDD GND NOR2_X1
xU11973 n912 n8287 n6420 VDD GND NOR2_X1
xU11974 n910 n8289 n6434 VDD GND NOR2_X1
xU11975 n909 n8288 n6441 VDD GND NOR2_X1
xU11976 n885 n8289 n6609 VDD GND NOR2_X1
xU11977 n892 n8288 n6560 VDD GND NOR2_X1
xU11978 n908 n8290 n6448 VDD GND NOR2_X1
xU11979 n905 n8290 n6469 VDD GND NOR2_X1
xU11980 n897 n8290 n6525 VDD GND NOR2_X1
xU11981 n891 n8290 n6567 VDD GND NOR2_X1
xU11982 n906 n8290 n6462 VDD GND NOR2_X1
xU11983 n900 n8290 n6504 VDD GND NOR2_X1
xU11984 n887 n8287 n6595 VDD GND NOR2_X1
xU11985 n907 n8290 n6455 VDD GND NOR2_X1
xU11986 n899 n8290 n6511 VDD GND NOR2_X1
xU11987 n890 n8286 n6574 VDD GND NOR2_X1
xU11988 n903 n8290 n6483 VDD GND NOR2_X1
xU11989 n896 n8290 n6532 VDD GND NOR2_X1
xU11990 n898 n8290 n6518 VDD GND NOR2_X1
xU11991 n888 n8289 n6588 VDD GND NOR2_X1
xU11992 n904 n8290 n6476 VDD GND NOR2_X1
xU11993 n895 n8288 n6539 VDD GND NOR2_X1
xU11994 n886 n8290 n6602 VDD GND NOR2_X1
xU11995 n902 n8290 n6490 VDD GND NOR2_X1
xU11996 n894 n8287 n6546 VDD GND NOR2_X1
xU11997 n889 n8286 n6581 VDD GND NOR2_X1
xU11998 n901 n8290 n6497 VDD GND NOR2_X1
xU11999 n893 n8289 n6553 VDD GND NOR2_X1
xU12000 n2669 n8347 n2667 VDD GND NOR2_X1
xU12001 n1651 n8349 n1649 VDD GND NOR2_X1
xU12002 n1420 n8350 n1418 VDD GND NOR2_X1
xU12003 n2474 n8348 n2472 VDD GND NOR2_X1
xU12004 n2240 n8348 n2238 VDD GND NOR2_X1
xU12005 n3489 n8346 n3487 VDD GND NOR2_X1
xU12006 n2645 n8347 n2643 VDD GND NOR2_X1
xU12007 n1442 n8350 n1440 VDD GND NOR2_X1
xU12008 n3536 n8346 n3534 VDD GND NOR2_X1
xU12009 n2844 n8346 n2842 VDD GND NOR2_X1
xU12010 n2898 n8346 n2896 VDD GND NOR2_X1
xU12011 n2289 n8348 n2287 VDD GND NOR2_X1
xU12012 n1228 n8350 n1226 VDD GND NOR2_X1
xU12013 n2991 n8346 n2989 VDD GND NOR2_X1
xU12014 n2265 n8348 n2263 VDD GND NOR2_X1
xU12015 n1204 n8350 n1202 VDD GND NOR2_X1
xU12016 n1397 n8350 n1395 VDD GND NOR2_X1
xU12017 n2523 n8348 n2521 VDD GND NOR2_X1
xU12018 n1275 n8350 n1273 VDD GND NOR2_X1
xU12019 n2453 n8348 n2451 VDD GND NOR2_X1
xU12020 n1743 n8349 n1741 VDD GND NOR2_X1
xU12021 n1327 n8350 n1325 VDD GND NOR2_X1
xU12022 n2572 n8347 n2570 VDD GND NOR2_X1
xU12023 n1354 n8350 n1352 VDD GND NOR2_X1
xU12024 n2546 n8347 n2544 VDD GND NOR2_X1
xU12025 n2695 n8347 n2693 VDD GND NOR2_X1
xU12026 n2775 n8347 n2773 VDD GND NOR2_X1
xU12027 n2802 n8347 n2800 VDD GND NOR2_X1
xU12028 n2726 n8347 n2724 VDD GND NOR2_X1
xU12029 n2822 n8347 n2820 VDD GND NOR2_X1
xU12030 n2372 n8348 n2370 VDD GND NOR2_X1
xU12031 n1621 n8349 n1619 VDD GND NOR2_X1
xU12032 n3562 n8346 n3560 VDD GND NOR2_X1
xU12033 n3514 n8346 n3512 VDD GND NOR2_X1
xU12034 n3108 n8346 n3106 VDD GND NOR2_X1
xU12035 n1596 n8349 n1594 VDD GND NOR2_X1
xU12036 n2498 n8348 n2496 VDD GND NOR2_X1
xU12037 n2751 n8347 n2749 VDD GND NOR2_X1
xU12038 n1807 n8349 n1805 VDD GND NOR2_X1
xU12039 n2869 n8346 n2867 VDD GND NOR2_X1
xU12040 n2429 n8348 n2427 VDD GND NOR2_X1
xU12041 n1722 n8349 n1720 VDD GND NOR2_X1
xU12042 n1472 n8350 n1470 VDD GND NOR2_X1
xU12043 n1524 n8349 n1522 VDD GND NOR2_X1
xU12044 n1552 n8349 n1550 VDD GND NOR2_X1
xU12045 n1574 n8349 n1572 VDD GND NOR2_X1
xU12046 n2970 n8346 n2968 VDD GND NOR2_X1
xU12047 n2216 n8349 n2214 VDD GND NOR2_X1
xU12048 n3053 n8346 n3051 VDD GND NOR2_X1
xU12049 n2344 n8348 n2342 VDD GND NOR2_X1
xU12050 n2317 n8348 n2315 VDD GND NOR2_X1
xU12051 n2403 n8348 n2401 VDD GND NOR2_X1
xU12052 n1373 n8350 n1371 VDD GND NOR2_X1
xU12053 n2600 n8347 n2598 VDD GND NOR2_X1
xU12054 n1302 n8350 n1300 VDD GND NOR2_X1
xU12055 n2622 n8347 n2620 VDD GND NOR2_X1
xU12056 n1249 n8350 n1247 VDD GND NOR2_X1
xU12057 n1495 n8349 n1493 VDD GND NOR2_X1
xU12058 n3463 n8346 n3461 VDD GND NOR2_X1
xU12059 n1862 n8349 n1860 VDD GND NOR2_X1
xU12060 n683 n8412 n7422 VDD GND NOR2_X1
xU12061 n684 n8412 n7392 VDD GND NOR2_X1
xU12062 n685 n8412 n7380 VDD GND NOR2_X1
xU12063 n785 n8422 n6102 VDD GND NOR2_X1
xU12064 n793 n8421 n6046 VDD GND NOR2_X1
xU12065 n761 n8419 n6270 VDD GND NOR2_X1
xU12066 n801 n8422 n5990 VDD GND NOR2_X1
xU12067 n769 n8420 n6214 VDD GND NOR2_X1
xU12068 n777 n8421 n6158 VDD GND NOR2_X1
xU12069 n781 n8421 n6130 VDD GND NOR2_X1
xU12070 n794 n8422 n6039 VDD GND NOR2_X1
xU12071 n762 n8419 n6263 VDD GND NOR2_X1
xU12072 n770 n8420 n6207 VDD GND NOR2_X1
xU12073 n778 n8421 n6151 VDD GND NOR2_X1
xU12074 n787 n8422 n6088 VDD GND NOR2_X1
xU12075 n796 n8422 n6025 VDD GND NOR2_X1
xU12076 n764 n8419 n6249 VDD GND NOR2_X1
xU12077 n773 n8420 n6186 VDD GND NOR2_X1
xU12078 n780 n8421 n6137 VDD GND NOR2_X1
xU12079 n788 n8420 n6081 VDD GND NOR2_X1
xU12080 n756 n8419 n6305 VDD GND NOR2_X1
xU12081 n795 n8422 n6032 VDD GND NOR2_X1
xU12082 n763 n8419 n6256 VDD GND NOR2_X1
xU12083 n776 n8421 n6165 VDD GND NOR2_X1
xU12084 n782 n8421 n6123 VDD GND NOR2_X1
xU12085 n791 n8420 n6060 VDD GND NOR2_X1
xU12086 n759 n8419 n6284 VDD GND NOR2_X1
xU12087 n799 n8422 n6004 VDD GND NOR2_X1
xU12088 n767 n8419 n6228 VDD GND NOR2_X1
xU12089 n803 n8421 n5976 VDD GND NOR2_X1
xU12090 n771 n8420 n6200 VDD GND NOR2_X1
xU12091 n779 n8420 n6144 VDD GND NOR2_X1
xU12092 n792 n8422 n6053 VDD GND NOR2_X1
xU12093 n760 n8419 n6277 VDD GND NOR2_X1
xU12094 n798 n8421 n6011 VDD GND NOR2_X1
xU12095 n766 n8419 n6235 VDD GND NOR2_X1
xU12096 n807 n8422 n5948 VDD GND NOR2_X1
xU12097 n775 n8421 n6172 VDD GND NOR2_X1
xU12098 n783 n8420 n6116 VDD GND NOR2_X1
xU12099 n789 n8422 n6074 VDD GND NOR2_X1
xU12100 n757 n8419 n6298 VDD GND NOR2_X1
xU12101 n800 n8422 n5997 VDD GND NOR2_X1
xU12102 n768 n8420 n6221 VDD GND NOR2_X1
xU12103 n774 n8420 n6179 VDD GND NOR2_X1
xU12104 n784 n8422 n6109 VDD GND NOR2_X1
xU12105 n797 n8421 n6018 VDD GND NOR2_X1
xU12106 n765 n8419 n6242 VDD GND NOR2_X1
xU12107 n790 n8420 n6067 VDD GND NOR2_X1
xU12108 n758 n8419 n6291 VDD GND NOR2_X1
xU12109 n804 n8421 n5969 VDD GND NOR2_X1
xU12110 n772 n8420 n6193 VDD GND NOR2_X1
xU12111 n802 n8423 n5983 VDD GND NOR2_X1
xU12112 n805 n8423 n5962 VDD GND NOR2_X1
xU12113 n808 n8423 n5939 VDD GND NOR2_X1
xU12114 n806 n8423 n5955 VDD GND NOR2_X1
xU12115 n7640 n7641 n8145 VDD GND NAND2_X1
xU12116 n8261 \AES_Comp_ENCa/Krg_32 n7640 VDD GND NAND2_X1
xU12117 n8279 Kin_32 n7641 VDD GND NAND2_X1
xU12118 n7638 n7639 n8144 VDD GND NAND2_X1
xU12119 n8261 \AES_Comp_ENCa/Krg_31 n7638 VDD GND NAND2_X1
xU12120 n8279 Kin_31 n7639 VDD GND NAND2_X1
xU12121 n7636 n7637 n8143 VDD GND NAND2_X1
xU12122 n8261 \AES_Comp_ENCa/Krg_30 n7636 VDD GND NAND2_X1
xU12123 n8279 Kin_30 n7637 VDD GND NAND2_X1
xU12124 n7634 n7635 n8142 VDD GND NAND2_X1
xU12125 n8261 \AES_Comp_ENCa/Krg_1 n7634 VDD GND NAND2_X1
xU12126 n8279 Kin_1 n7635 VDD GND NAND2_X1
xU12127 n7632 n7633 n8141 VDD GND NAND2_X1
xU12128 n8260 \AES_Comp_ENCa/Krg_29 n7632 VDD GND NAND2_X1
xU12129 n8279 Kin_29 n7633 VDD GND NAND2_X1
xU12130 n7630 n7631 n8140 VDD GND NAND2_X1
xU12131 n8260 \AES_Comp_ENCa/Krg_28 n7630 VDD GND NAND2_X1
xU12132 n8279 Kin_28 n7631 VDD GND NAND2_X1
xU12133 n7628 n7629 n8139 VDD GND NAND2_X1
xU12134 n8260 \AES_Comp_ENCa/Krg_27 n7628 VDD GND NAND2_X1
xU12135 n8279 Kin_27 n7629 VDD GND NAND2_X1
xU12136 n7626 n7627 n8138 VDD GND NAND2_X1
xU12137 n8260 \AES_Comp_ENCa/Krg_26 n7626 VDD GND NAND2_X1
xU12138 n8279 Kin_26 n7627 VDD GND NAND2_X1
xU12139 n7624 n7625 n8137 VDD GND NAND2_X1
xU12140 n8260 \AES_Comp_ENCa/Krg_25 n7624 VDD GND NAND2_X1
xU12141 n8279 Kin_25 n7625 VDD GND NAND2_X1
xU12142 n7622 n7623 n8136 VDD GND NAND2_X1
xU12143 n8260 \AES_Comp_ENCa/Krg_24 n7622 VDD GND NAND2_X1
xU12144 n8279 Kin_24 n7623 VDD GND NAND2_X1
xU12145 n7620 n7621 n8135 VDD GND NAND2_X1
xU12146 n8260 \AES_Comp_ENCa/Krg_23 n7620 VDD GND NAND2_X1
xU12147 n8279 Kin_23 n7621 VDD GND NAND2_X1
xU12148 n7618 n7619 n8134 VDD GND NAND2_X1
xU12149 n8260 \AES_Comp_ENCa/Krg_22 n7618 VDD GND NAND2_X1
xU12150 n8279 Kin_22 n7619 VDD GND NAND2_X1
xU12151 n7616 n7617 n8133 VDD GND NAND2_X1
xU12152 n8260 \AES_Comp_ENCa/Krg_21 n7616 VDD GND NAND2_X1
xU12153 n8280 Kin_21 n7617 VDD GND NAND2_X1
xU12154 n7614 n7615 n8132 VDD GND NAND2_X1
xU12155 n8260 \AES_Comp_ENCa/Krg_20 n7614 VDD GND NAND2_X1
xU12156 n8280 Kin_20 n7615 VDD GND NAND2_X1
xU12157 n7612 n7613 n8131 VDD GND NAND2_X1
xU12158 n8259 \AES_Comp_ENCa/Krg_19 n7612 VDD GND NAND2_X1
xU12159 n8280 Kin_19 n7613 VDD GND NAND2_X1
xU12160 n7610 n7611 n8130 VDD GND NAND2_X1
xU12161 n8259 \AES_Comp_ENCa/Krg_18 n7610 VDD GND NAND2_X1
xU12162 n8280 Kin_18 n7611 VDD GND NAND2_X1
xU12163 n7608 n7609 n8129 VDD GND NAND2_X1
xU12164 n8259 \AES_Comp_ENCa/Krg_17 n7608 VDD GND NAND2_X1
xU12165 n8280 Kin_17 n7609 VDD GND NAND2_X1
xU12166 n7606 n7607 n8128 VDD GND NAND2_X1
xU12167 n8259 \AES_Comp_ENCa/Krg_16 n7606 VDD GND NAND2_X1
xU12168 n8280 Kin_16 n7607 VDD GND NAND2_X1
xU12169 n7604 n7605 n8127 VDD GND NAND2_X1
xU12170 n8259 \AES_Comp_ENCa/Krg_15 n7604 VDD GND NAND2_X1
xU12171 n8280 Kin_15 n7605 VDD GND NAND2_X1
xU12172 n7602 n7603 n8126 VDD GND NAND2_X1
xU12173 n8259 \AES_Comp_ENCa/Krg_14 n7602 VDD GND NAND2_X1
xU12174 n8280 Kin_14 n7603 VDD GND NAND2_X1
xU12175 n7600 n7601 n8125 VDD GND NAND2_X1
xU12176 n8259 \AES_Comp_ENCa/Krg_13 n7600 VDD GND NAND2_X1
xU12177 n8280 Kin_13 n7601 VDD GND NAND2_X1
xU12178 n7598 n7599 n8124 VDD GND NAND2_X1
xU12179 n8259 \AES_Comp_ENCa/Krg_12 n7598 VDD GND NAND2_X1
xU12180 n8280 Kin_12 n7599 VDD GND NAND2_X1
xU12181 n7596 n7597 n8123 VDD GND NAND2_X1
xU12182 n8259 \AES_Comp_ENCa/Krg_11 n7596 VDD GND NAND2_X1
xU12183 n8280 Kin_11 n7597 VDD GND NAND2_X1
xU12184 n7594 n7595 n8122 VDD GND NAND2_X1
xU12185 n8259 \AES_Comp_ENCa/Krg_10 n7594 VDD GND NAND2_X1
xU12186 n8280 Kin_10 n7595 VDD GND NAND2_X1
xU12187 n7835 n7836 n8243 VDD GND NAND2_X1
xU12188 n8258 \AES_Comp_ENCa/Krg_0 n7835 VDD GND NAND2_X1
xU12189 n8272 Kin_0 n7836 VDD GND NAND2_X1
xU12190 n7830 n7831 n8240 VDD GND NAND2_X1
xU12191 n8270 \AES_Comp_ENCa/Krg_127 n7830 VDD GND NAND2_X1
xU12192 n8272 Kin_127 n7831 VDD GND NAND2_X1
xU12193 n7828 n7829 n8239 VDD GND NAND2_X1
xU12194 n8270 \AES_Comp_ENCa/Krg_126 n7828 VDD GND NAND2_X1
xU12195 n8272 Kin_126 n7829 VDD GND NAND2_X1
xU12196 n7826 n7827 n8238 VDD GND NAND2_X1
xU12197 n8270 \AES_Comp_ENCa/Krg_125 n7826 VDD GND NAND2_X1
xU12198 n8272 Kin_125 n7827 VDD GND NAND2_X1
xU12199 n7824 n7825 n8237 VDD GND NAND2_X1
xU12200 n8270 \AES_Comp_ENCa/Krg_124 n7824 VDD GND NAND2_X1
xU12201 n8272 Kin_124 n7825 VDD GND NAND2_X1
xU12202 n7822 n7823 n8236 VDD GND NAND2_X1
xU12203 n8270 \AES_Comp_ENCa/Krg_123 n7822 VDD GND NAND2_X1
xU12204 n8272 Kin_123 n7823 VDD GND NAND2_X1
xU12205 n7820 n7821 n8235 VDD GND NAND2_X1
xU12206 n8270 \AES_Comp_ENCa/Krg_122 n7820 VDD GND NAND2_X1
xU12207 n8272 Kin_122 n7821 VDD GND NAND2_X1
xU12208 n7818 n7819 n8234 VDD GND NAND2_X1
xU12209 n8270 \AES_Comp_ENCa/Krg_121 n7818 VDD GND NAND2_X1
xU12210 n8272 Kin_121 n7819 VDD GND NAND2_X1
xU12211 n7816 n7817 n8233 VDD GND NAND2_X1
xU12212 n8270 \AES_Comp_ENCa/Krg_120 n7816 VDD GND NAND2_X1
xU12213 n8272 Kin_120 n7817 VDD GND NAND2_X1
xU12214 n7814 n7815 n8232 VDD GND NAND2_X1
xU12215 n8270 \AES_Comp_ENCa/Krg_119 n7814 VDD GND NAND2_X1
xU12216 n8272 Kin_119 n7815 VDD GND NAND2_X1
xU12217 n7812 n7813 n8231 VDD GND NAND2_X1
xU12218 n8270 \AES_Comp_ENCa/Krg_118 n7812 VDD GND NAND2_X1
xU12219 n8272 Kin_118 n7813 VDD GND NAND2_X1
xU12220 n7810 n7811 n8230 VDD GND NAND2_X1
xU12221 n8269 \AES_Comp_ENCa/Krg_117 n7810 VDD GND NAND2_X1
xU12222 n8272 Kin_117 n7811 VDD GND NAND2_X1
xU12223 n7808 n7809 n8229 VDD GND NAND2_X1
xU12224 n8269 \AES_Comp_ENCa/Krg_116 n7808 VDD GND NAND2_X1
xU12225 n8273 Kin_116 n7809 VDD GND NAND2_X1
xU12226 n7806 n7807 n8228 VDD GND NAND2_X1
xU12227 n8269 \AES_Comp_ENCa/Krg_115 n7806 VDD GND NAND2_X1
xU12228 n8273 Kin_115 n7807 VDD GND NAND2_X1
xU12229 n7804 n7805 n8227 VDD GND NAND2_X1
xU12230 n8269 \AES_Comp_ENCa/Krg_114 n7804 VDD GND NAND2_X1
xU12231 n8273 Kin_114 n7805 VDD GND NAND2_X1
xU12232 n7802 n7803 n8226 VDD GND NAND2_X1
xU12233 n8269 \AES_Comp_ENCa/Krg_113 n7802 VDD GND NAND2_X1
xU12234 n8273 Kin_113 n7803 VDD GND NAND2_X1
xU12235 n7800 n7801 n8225 VDD GND NAND2_X1
xU12236 n8269 \AES_Comp_ENCa/Krg_112 n7800 VDD GND NAND2_X1
xU12237 n8273 Kin_112 n7801 VDD GND NAND2_X1
xU12238 n7798 n7799 n8224 VDD GND NAND2_X1
xU12239 n8269 \AES_Comp_ENCa/Krg_111 n7798 VDD GND NAND2_X1
xU12240 n8273 Kin_111 n7799 VDD GND NAND2_X1
xU12241 n7796 n7797 n8223 VDD GND NAND2_X1
xU12242 n8269 \AES_Comp_ENCa/Krg_110 n7796 VDD GND NAND2_X1
xU12243 n8273 Kin_110 n7797 VDD GND NAND2_X1
xU12244 n7794 n7795 n8222 VDD GND NAND2_X1
xU12245 n8269 \AES_Comp_ENCa/Krg_109 n7794 VDD GND NAND2_X1
xU12246 n8273 Kin_109 n7795 VDD GND NAND2_X1
xU12247 n7792 n7793 n8221 VDD GND NAND2_X1
xU12248 n8269 \AES_Comp_ENCa/Krg_108 n7792 VDD GND NAND2_X1
xU12249 n8273 Kin_108 n7793 VDD GND NAND2_X1
xU12250 n7790 n7791 n8220 VDD GND NAND2_X1
xU12251 n8268 \AES_Comp_ENCa/Krg_107 n7790 VDD GND NAND2_X1
xU12252 n8273 Kin_107 n7791 VDD GND NAND2_X1
xU12253 n7788 n7789 n8219 VDD GND NAND2_X1
xU12254 n8268 \AES_Comp_ENCa/Krg_106 n7788 VDD GND NAND2_X1
xU12255 n8273 Kin_106 n7789 VDD GND NAND2_X1
xU12256 n7786 n7787 n8218 VDD GND NAND2_X1
xU12257 n8268 \AES_Comp_ENCa/Krg_105 n7786 VDD GND NAND2_X1
xU12258 n8273 Kin_105 n7787 VDD GND NAND2_X1
xU12259 n7784 n7785 n8217 VDD GND NAND2_X1
xU12260 n8268 \AES_Comp_ENCa/Krg_104 n7784 VDD GND NAND2_X1
xU12261 n8274 Kin_104 n7785 VDD GND NAND2_X1
xU12262 n7782 n7783 n8216 VDD GND NAND2_X1
xU12263 n8268 \AES_Comp_ENCa/Krg_103 n7782 VDD GND NAND2_X1
xU12264 n8274 Kin_103 n7783 VDD GND NAND2_X1
xU12265 n7780 n7781 n8215 VDD GND NAND2_X1
xU12266 n8268 \AES_Comp_ENCa/Krg_102 n7780 VDD GND NAND2_X1
xU12267 n8274 Kin_102 n7781 VDD GND NAND2_X1
xU12268 n7778 n7779 n8214 VDD GND NAND2_X1
xU12269 n8268 \AES_Comp_ENCa/Krg_101 n7778 VDD GND NAND2_X1
xU12270 n8274 Kin_101 n7779 VDD GND NAND2_X1
xU12271 n7776 n7777 n8213 VDD GND NAND2_X1
xU12272 n8268 \AES_Comp_ENCa/Krg_100 n7776 VDD GND NAND2_X1
xU12273 n8274 Kin_100 n7777 VDD GND NAND2_X1
xU12274 n7774 n7775 n8212 VDD GND NAND2_X1
xU12275 n8268 \AES_Comp_ENCa/Krg_99 n7774 VDD GND NAND2_X1
xU12276 n8274 Kin_99 n7775 VDD GND NAND2_X1
xU12277 n7772 n7773 n8211 VDD GND NAND2_X1
xU12278 n8268 \AES_Comp_ENCa/Krg_98 n7772 VDD GND NAND2_X1
xU12279 n8274 Kin_98 n7773 VDD GND NAND2_X1
xU12280 n7770 n7771 n8210 VDD GND NAND2_X1
xU12281 n8267 \AES_Comp_ENCa/Krg_97 n7770 VDD GND NAND2_X1
xU12282 n8274 Kin_97 n7771 VDD GND NAND2_X1
xU12283 n7768 n7769 n8209 VDD GND NAND2_X1
xU12284 n8267 \AES_Comp_ENCa/Krg_96 n7768 VDD GND NAND2_X1
xU12285 n8274 Kin_96 n7769 VDD GND NAND2_X1
xU12286 n7766 n7767 n8208 VDD GND NAND2_X1
xU12287 n8267 \AES_Comp_ENCa/Krg_95 n7766 VDD GND NAND2_X1
xU12288 n8274 Kin_95 n7767 VDD GND NAND2_X1
xU12289 n7764 n7765 n8207 VDD GND NAND2_X1
xU12290 n8267 \AES_Comp_ENCa/Krg_94 n7764 VDD GND NAND2_X1
xU12291 n8274 Kin_94 n7765 VDD GND NAND2_X1
xU12292 n7762 n7763 n8206 VDD GND NAND2_X1
xU12293 n8267 \AES_Comp_ENCa/Krg_93 n7762 VDD GND NAND2_X1
xU12294 n8274 Kin_93 n7763 VDD GND NAND2_X1
xU12295 n7760 n7761 n8205 VDD GND NAND2_X1
xU12296 n8267 \AES_Comp_ENCa/Krg_92 n7760 VDD GND NAND2_X1
xU12297 n8275 Kin_92 n7761 VDD GND NAND2_X1
xU12298 n7758 n7759 n8204 VDD GND NAND2_X1
xU12299 n8267 \AES_Comp_ENCa/Krg_91 n7758 VDD GND NAND2_X1
xU12300 n8275 Kin_91 n7759 VDD GND NAND2_X1
xU12301 n7756 n7757 n8203 VDD GND NAND2_X1
xU12302 n8267 \AES_Comp_ENCa/Krg_90 n7756 VDD GND NAND2_X1
xU12303 n8275 Kin_90 n7757 VDD GND NAND2_X1
xU12304 n7754 n7755 n8202 VDD GND NAND2_X1
xU12305 n8267 \AES_Comp_ENCa/Krg_89 n7754 VDD GND NAND2_X1
xU12306 n8275 Kin_89 n7755 VDD GND NAND2_X1
xU12307 n7752 n7753 n8201 VDD GND NAND2_X1
xU12308 n8267 \AES_Comp_ENCa/Krg_88 n7752 VDD GND NAND2_X1
xU12309 n8275 Kin_88 n7753 VDD GND NAND2_X1
xU12310 n7750 n7751 n8200 VDD GND NAND2_X1
xU12311 n8266 \AES_Comp_ENCa/Krg_87 n7750 VDD GND NAND2_X1
xU12312 n8275 Kin_87 n7751 VDD GND NAND2_X1
xU12313 n7748 n7749 n8199 VDD GND NAND2_X1
xU12314 n8266 \AES_Comp_ENCa/Krg_86 n7748 VDD GND NAND2_X1
xU12315 n8275 Kin_86 n7749 VDD GND NAND2_X1
xU12316 n7746 n7747 n8198 VDD GND NAND2_X1
xU12317 n8266 \AES_Comp_ENCa/Krg_85 n7746 VDD GND NAND2_X1
xU12318 n8275 Kin_85 n7747 VDD GND NAND2_X1
xU12319 n7744 n7745 n8197 VDD GND NAND2_X1
xU12320 n8266 \AES_Comp_ENCa/Krg_84 n7744 VDD GND NAND2_X1
xU12321 n8275 Kin_84 n7745 VDD GND NAND2_X1
xU12322 n7742 n7743 n8196 VDD GND NAND2_X1
xU12323 n8266 \AES_Comp_ENCa/Krg_83 n7742 VDD GND NAND2_X1
xU12324 n8275 Kin_83 n7743 VDD GND NAND2_X1
xU12325 n7740 n7741 n8195 VDD GND NAND2_X1
xU12326 n8266 \AES_Comp_ENCa/Krg_82 n7740 VDD GND NAND2_X1
xU12327 n8275 Kin_82 n7741 VDD GND NAND2_X1
xU12328 n7738 n7739 n8194 VDD GND NAND2_X1
xU12329 n8266 \AES_Comp_ENCa/Krg_81 n7738 VDD GND NAND2_X1
xU12330 n8275 Kin_81 n7739 VDD GND NAND2_X1
xU12331 n7736 n7737 n8193 VDD GND NAND2_X1
xU12332 n8266 \AES_Comp_ENCa/Krg_80 n7736 VDD GND NAND2_X1
xU12333 n8276 Kin_80 n7737 VDD GND NAND2_X1
xU12334 n7734 n7735 n8192 VDD GND NAND2_X1
xU12335 n8266 \AES_Comp_ENCa/Krg_79 n7734 VDD GND NAND2_X1
xU12336 n8276 Kin_79 n7735 VDD GND NAND2_X1
xU12337 n7732 n7733 n8191 VDD GND NAND2_X1
xU12338 n8266 \AES_Comp_ENCa/Krg_78 n7732 VDD GND NAND2_X1
xU12339 n8276 Kin_78 n7733 VDD GND NAND2_X1
xU12340 n7730 n7731 n8190 VDD GND NAND2_X1
xU12341 n8265 \AES_Comp_ENCa/Krg_77 n7730 VDD GND NAND2_X1
xU12342 n8276 Kin_77 n7731 VDD GND NAND2_X1
xU12343 n7728 n7729 n8189 VDD GND NAND2_X1
xU12344 n8265 \AES_Comp_ENCa/Krg_76 n7728 VDD GND NAND2_X1
xU12345 n8276 Kin_76 n7729 VDD GND NAND2_X1
xU12346 n7726 n7727 n8188 VDD GND NAND2_X1
xU12347 n8265 \AES_Comp_ENCa/Krg_75 n7726 VDD GND NAND2_X1
xU12348 n8276 Kin_75 n7727 VDD GND NAND2_X1
xU12349 n7724 n7725 n8187 VDD GND NAND2_X1
xU12350 n8265 \AES_Comp_ENCa/Krg_74 n7724 VDD GND NAND2_X1
xU12351 n8276 Kin_74 n7725 VDD GND NAND2_X1
xU12352 n7722 n7723 n8186 VDD GND NAND2_X1
xU12353 n8265 \AES_Comp_ENCa/Krg_73 n7722 VDD GND NAND2_X1
xU12354 n8276 Kin_73 n7723 VDD GND NAND2_X1
xU12355 n7720 n7721 n8185 VDD GND NAND2_X1
xU12356 n8265 \AES_Comp_ENCa/Krg_72 n7720 VDD GND NAND2_X1
xU12357 n8276 Kin_72 n7721 VDD GND NAND2_X1
xU12358 n7718 n7719 n8184 VDD GND NAND2_X1
xU12359 n8265 \AES_Comp_ENCa/Krg_71 n7718 VDD GND NAND2_X1
xU12360 n8276 Kin_71 n7719 VDD GND NAND2_X1
xU12361 n7716 n7717 n8183 VDD GND NAND2_X1
xU12362 n8265 \AES_Comp_ENCa/Krg_70 n7716 VDD GND NAND2_X1
xU12363 n8276 Kin_70 n7717 VDD GND NAND2_X1
xU12364 n7714 n7715 n8182 VDD GND NAND2_X1
xU12365 n8265 \AES_Comp_ENCa/Krg_69 n7714 VDD GND NAND2_X1
xU12366 n8276 Kin_69 n7715 VDD GND NAND2_X1
xU12367 n7712 n7713 n8181 VDD GND NAND2_X1
xU12368 n8265 \AES_Comp_ENCa/Krg_68 n7712 VDD GND NAND2_X1
xU12369 n8277 Kin_68 n7713 VDD GND NAND2_X1
xU12370 n7710 n7711 n8180 VDD GND NAND2_X1
xU12371 n8264 \AES_Comp_ENCa/Krg_67 n7710 VDD GND NAND2_X1
xU12372 n8277 Kin_67 n7711 VDD GND NAND2_X1
xU12373 n7708 n7709 n8179 VDD GND NAND2_X1
xU12374 n8264 \AES_Comp_ENCa/Krg_66 n7708 VDD GND NAND2_X1
xU12375 n8277 Kin_66 n7709 VDD GND NAND2_X1
xU12376 n7706 n7707 n8178 VDD GND NAND2_X1
xU12377 n8264 \AES_Comp_ENCa/Krg_65 n7706 VDD GND NAND2_X1
xU12378 n8277 Kin_65 n7707 VDD GND NAND2_X1
xU12379 n7704 n7705 n8177 VDD GND NAND2_X1
xU12380 n8264 \AES_Comp_ENCa/Krg_64 n7704 VDD GND NAND2_X1
xU12381 n8277 Kin_64 n7705 VDD GND NAND2_X1
xU12382 n7702 n7703 n8176 VDD GND NAND2_X1
xU12383 n8264 \AES_Comp_ENCa/Krg_63 n7702 VDD GND NAND2_X1
xU12384 n8277 Kin_63 n7703 VDD GND NAND2_X1
xU12385 n7700 n7701 n8175 VDD GND NAND2_X1
xU12386 n8264 \AES_Comp_ENCa/Krg_62 n7700 VDD GND NAND2_X1
xU12387 n8277 Kin_62 n7701 VDD GND NAND2_X1
xU12388 n7698 n7699 n8174 VDD GND NAND2_X1
xU12389 n8264 \AES_Comp_ENCa/Krg_61 n7698 VDD GND NAND2_X1
xU12390 n8277 Kin_61 n7699 VDD GND NAND2_X1
xU12391 n7696 n7697 n8173 VDD GND NAND2_X1
xU12392 n8264 \AES_Comp_ENCa/Krg_60 n7696 VDD GND NAND2_X1
xU12393 n8277 Kin_60 n7697 VDD GND NAND2_X1
xU12394 n7694 n7695 n8172 VDD GND NAND2_X1
xU12395 n8264 \AES_Comp_ENCa/Krg_59 n7694 VDD GND NAND2_X1
xU12396 n8277 Kin_59 n7695 VDD GND NAND2_X1
xU12397 n7692 n7693 n8171 VDD GND NAND2_X1
xU12398 n8263 \AES_Comp_ENCa/Krg_58 n7692 VDD GND NAND2_X1
xU12399 n8277 Kin_58 n7693 VDD GND NAND2_X1
xU12400 n7690 n7691 n8170 VDD GND NAND2_X1
xU12401 n8263 \AES_Comp_ENCa/Krg_57 n7690 VDD GND NAND2_X1
xU12402 n8277 Kin_57 n7691 VDD GND NAND2_X1
xU12403 n7688 n7689 n8169 VDD GND NAND2_X1
xU12404 n8263 \AES_Comp_ENCa/Krg_56 n7688 VDD GND NAND2_X1
xU12405 n8278 Kin_56 n7689 VDD GND NAND2_X1
xU12406 n7686 n7687 n8168 VDD GND NAND2_X1
xU12407 n8263 \AES_Comp_ENCa/Krg_55 n7686 VDD GND NAND2_X1
xU12408 n8278 Kin_55 n7687 VDD GND NAND2_X1
xU12409 n7684 n7685 n8167 VDD GND NAND2_X1
xU12410 n8263 \AES_Comp_ENCa/Krg_54 n7684 VDD GND NAND2_X1
xU12411 n8278 Kin_54 n7685 VDD GND NAND2_X1
xU12412 n7682 n7683 n8166 VDD GND NAND2_X1
xU12413 n8263 \AES_Comp_ENCa/Krg_53 n7682 VDD GND NAND2_X1
xU12414 n8278 Kin_53 n7683 VDD GND NAND2_X1
xU12415 n7680 n7681 n8165 VDD GND NAND2_X1
xU12416 n8263 \AES_Comp_ENCa/Krg_52 n7680 VDD GND NAND2_X1
xU12417 n8278 Kin_52 n7681 VDD GND NAND2_X1
xU12418 n7678 n7679 n8164 VDD GND NAND2_X1
xU12419 n8263 \AES_Comp_ENCa/Krg_51 n7678 VDD GND NAND2_X1
xU12420 n8278 Kin_51 n7679 VDD GND NAND2_X1
xU12421 n7676 n7677 n8163 VDD GND NAND2_X1
xU12422 n8263 \AES_Comp_ENCa/Krg_50 n7676 VDD GND NAND2_X1
xU12423 n8278 Kin_50 n7677 VDD GND NAND2_X1
xU12424 n7674 n7675 n8162 VDD GND NAND2_X1
xU12425 n8263 \AES_Comp_ENCa/Krg_49 n7674 VDD GND NAND2_X1
xU12426 n8278 Kin_49 n7675 VDD GND NAND2_X1
xU12427 n7672 n7673 n8161 VDD GND NAND2_X1
xU12428 n8262 \AES_Comp_ENCa/Krg_48 n7672 VDD GND NAND2_X1
xU12429 n8278 Kin_48 n7673 VDD GND NAND2_X1
xU12430 n7670 n7671 n8160 VDD GND NAND2_X1
xU12431 n8262 \AES_Comp_ENCa/Krg_47 n7670 VDD GND NAND2_X1
xU12432 n8278 Kin_47 n7671 VDD GND NAND2_X1
xU12433 n7668 n7669 n8159 VDD GND NAND2_X1
xU12434 n8262 \AES_Comp_ENCa/Krg_46 n7668 VDD GND NAND2_X1
xU12435 n8278 Kin_46 n7669 VDD GND NAND2_X1
xU12436 n7666 n7667 n8158 VDD GND NAND2_X1
xU12437 n8262 \AES_Comp_ENCa/Krg_45 n7666 VDD GND NAND2_X1
xU12438 n8278 Kin_45 n7667 VDD GND NAND2_X1
xU12439 n7664 n7665 n8157 VDD GND NAND2_X1
xU12440 n8262 \AES_Comp_ENCa/Krg_44 n7664 VDD GND NAND2_X1
xU12441 n7578 Kin_44 n7665 VDD GND NAND2_X1
xU12442 n7662 n7663 n8156 VDD GND NAND2_X1
xU12443 n8262 \AES_Comp_ENCa/Krg_43 n7662 VDD GND NAND2_X1
xU12444 n8271 Kin_43 n7663 VDD GND NAND2_X1
xU12445 n7660 n7661 n8155 VDD GND NAND2_X1
xU12446 n8262 \AES_Comp_ENCa/Krg_42 n7660 VDD GND NAND2_X1
xU12447 n7578 Kin_42 n7661 VDD GND NAND2_X1
xU12448 n7658 n7659 n8154 VDD GND NAND2_X1
xU12449 n8262 \AES_Comp_ENCa/Krg_41 n7658 VDD GND NAND2_X1
xU12450 n8271 Kin_41 n7659 VDD GND NAND2_X1
xU12451 n7656 n7657 n8153 VDD GND NAND2_X1
xU12452 n8262 \AES_Comp_ENCa/Krg_40 n7656 VDD GND NAND2_X1
xU12453 n7578 Kin_40 n7657 VDD GND NAND2_X1
xU12454 n7654 n7655 n8152 VDD GND NAND2_X1
xU12455 n8262 \AES_Comp_ENCa/Krg_39 n7654 VDD GND NAND2_X1
xU12456 n7578 Kin_39 n7655 VDD GND NAND2_X1
xU12457 n7652 n7653 n8151 VDD GND NAND2_X1
xU12458 n8261 \AES_Comp_ENCa/Krg_38 n7652 VDD GND NAND2_X1
xU12459 n7578 Kin_38 n7653 VDD GND NAND2_X1
xU12460 n7650 n7651 n8150 VDD GND NAND2_X1
xU12461 n8261 \AES_Comp_ENCa/Krg_37 n7650 VDD GND NAND2_X1
xU12462 n7578 Kin_37 n7651 VDD GND NAND2_X1
xU12463 n7648 n7649 n8149 VDD GND NAND2_X1
xU12464 n8261 \AES_Comp_ENCa/Krg_36 n7648 VDD GND NAND2_X1
xU12465 n8271 Kin_36 n7649 VDD GND NAND2_X1
xU12466 n7646 n7647 n8148 VDD GND NAND2_X1
xU12467 n8261 \AES_Comp_ENCa/Krg_35 n7646 VDD GND NAND2_X1
xU12468 n8271 Kin_35 n7647 VDD GND NAND2_X1
xU12469 n7644 n7645 n8147 VDD GND NAND2_X1
xU12470 n8261 \AES_Comp_ENCa/Krg_34 n7644 VDD GND NAND2_X1
xU12471 n8271 Kin_34 n7645 VDD GND NAND2_X1
xU12472 n7642 n7643 n8146 VDD GND NAND2_X1
xU12473 n8261 \AES_Comp_ENCa/Krg_33 n7642 VDD GND NAND2_X1
xU12474 n8271 Kin_33 n7643 VDD GND NAND2_X1
xU12475 \AES_Comp_ENCa/Rrg_1 n813 n6766 VDD GND NAND2_X1
xU12476 Krdy n5935 n5944 VDD GND NAND2_X1
xU12477 n7453 RSTn n1007 VDD GND NAND2_X1
xU12478 n5931 n7454 n7453 VDD GND NOR2_X1
xU12479 n7452 n7455 n7454 VDD GND NOR2_X1
xU12480 n7564 n7565 n8111 VDD GND NAND2_X1
xU12481 n7566 n809 n7564 VDD GND OR2_X1
xU12482 n5931 n7566 n7565 VDD GND NAND2_X1
xU12483 n130 n8313 n7566 VDD GND NAND2_X1
xU12484 RSTn n8325 n7579 VDD GND AND2_X1
xU12485 n7832 n7833 n8241 VDD GND NAND2_X1
xU12486 Kvld_reg n7563 n7832 VDD GND NAND2_X1
xU12487 Kvld_E n136 n7833 VDD GND NAND2_X1
xU12488 n7840 RSTn n7839 VDD GND NAND2_X1
xU12489 n7841 n7842 n7840 VDD GND NOR2_X1
xU12490 n133 n5935 n7842 VDD GND AND2_X1
xU12491 n5931 \AES_Comp_ENCa/Rrg_0 n7841 VDD GND AND2_X1
xU12492 n8281 n7834 n8242 VDD GND NAND2_X1
xU12493 Kvld_E n8258 n7834 VDD GND NAND2_X1
xU12494 n7592 n7593 n8121 VDD GND NAND2_X1
xU12495 n8258 \AES_Comp_ENCa/Krg_9 n7592 VDD GND NAND2_X1
xU12496 n8271 Kin_9 n7593 VDD GND NAND2_X1
xU12497 n7590 n7591 n8120 VDD GND NAND2_X1
xU12498 n8258 \AES_Comp_ENCa/Krg_8 n7590 VDD GND NAND2_X1
xU12499 n7578 Kin_8 n7591 VDD GND NAND2_X1
xU12500 n7588 n7589 n8119 VDD GND NAND2_X1
xU12501 n8258 \AES_Comp_ENCa/Krg_7 n7588 VDD GND NAND2_X1
xU12502 n7578 Kin_7 n7589 VDD GND NAND2_X1
xU12503 n7586 n7587 n8118 VDD GND NAND2_X1
xU12504 n8258 \AES_Comp_ENCa/Krg_6 n7586 VDD GND NAND2_X1
xU12505 n8271 Kin_6 n7587 VDD GND NAND2_X1
xU12506 n7584 n7585 n8117 VDD GND NAND2_X1
xU12507 n8258 \AES_Comp_ENCa/Krg_5 n7584 VDD GND NAND2_X1
xU12508 n7578 Kin_5 n7585 VDD GND NAND2_X1
xU12509 n7582 n7583 n8116 VDD GND NAND2_X1
xU12510 n8258 \AES_Comp_ENCa/Krg_4 n7582 VDD GND NAND2_X1
xU12511 n8271 Kin_4 n7583 VDD GND NAND2_X1
xU12512 n7580 n7581 n8115 VDD GND NAND2_X1
xU12513 n8258 \AES_Comp_ENCa/Krg_3 n7580 VDD GND NAND2_X1
xU12514 n7578 Kin_3 n7581 VDD GND NAND2_X1
xU12515 n7576 n7577 n8114 VDD GND NAND2_X1
xU12516 n8264 \AES_Comp_ENCa/Krg_2 n7576 VDD GND NAND2_X1
xU12517 n8271 Kin_2 n7577 VDD GND NAND2_X1
xU12518 n7837 n7838 n8244 VDD GND NAND2_X1
xU12519 n5935 n7839 n7838 VDD GND NAND2_X1
xU12520 n130 BSY_E n7837 VDD GND NAND2_X1
xU12521 n7561 n7562 n8110 VDD GND NAND2_X1
xU12522 Dvld_reg n7563 n7561 VDD GND NAND2_X1
xU12523 Dvld_E n136 n7562 VDD GND NAND2_X1
xU12524 n7843 RSTn n7452 VDD GND NAND2_X1
xU12525 n8434 n137 n7843 VDD GND NOR2_X1
xU12526 EncDec n8437 VDD GND BUF_X1
xU12527 EncDec n8438 VDD GND BUF_X1
xU12528 EncDec n8439 VDD GND BUF_X1
xU12529 EncDec n8440 VDD GND BUF_X1
xU12530 EncDec n8441 VDD GND BUF_X1
xU12531 EncDec n8442 VDD GND BUF_X1
xU12532 EncDec n8443 VDD GND BUF_X1
xU12533 EncDec n8434 VDD GND BUF_X1
xU12534 EncDec n8435 VDD GND BUF_X1
xU12535 EncDec n8436 VDD GND BUF_X1
xU12536 EncDec n8444 VDD GND BUF_X1
xU12537 Drdy n135 n7455 VDD GND NAND2_X1
xU12538 RSTn n137 n7563 VDD GND AND2_X1
xU12539 n8437 n362 Dout_25 VDD GND NOR2_X1
xU12540 n8444 n593 Dout_97 VDD GND NOR2_X1
xU12541 n8438 n367 Dout_29 VDD GND NOR2_X1
xU12542 n8434 n618 Dout_105 VDD GND NOR2_X1
xU12543 Krdy n135 VDD GND INV_X1
xU12544 n8437 n190 Dout_1 VDD GND NOR2_X1
xU12545 n8442 n520 Dout_79 VDD GND NOR2_X1
xU12546 n8441 n485 Dout_65 VDD GND NOR2_X1
xU12547 n8435 n653 Dout_116 VDD GND NOR2_X1
xU12548 n8440 n434 Dout_49 VDD GND NOR2_X1
xU12549 n8444 n245 Dout_9 VDD GND NOR2_X1
xU12550 n8443 n243 Dout_8 VDD GND NOR2_X1
xU12551 n8444 n591 Dout_96 VDD GND NOR2_X1
xU12552 n8440 n194 Dout_4 VDD GND NOR2_X1
xU12553 n8436 n677 Dout_124 VDD GND NOR2_X1
xU12554 n8436 n680 Dout_127 VDD GND NOR2_X1
xU12555 n8436 n255 Dout_15 VDD GND NOR2_X1
xU12556 n8438 n366 Dout_28 VDD GND NOR2_X1
xU12557 n8438 n392 Dout_36 VDD GND NOR2_X1
xU12558 n8440 n440 Dout_52 VDD GND NOR2_X1
xU12559 n8441 n465 Dout_60 VDD GND NOR2_X1
xU12560 n8441 n468 Dout_63 VDD GND NOR2_X1
xU12561 n8441 n492 Dout_68 VDD GND NOR2_X1
xU12562 n8442 n517 Dout_76 VDD GND NOR2_X1
xU12563 n8444 n568 Dout_92 VDD GND NOR2_X1
xU12564 n8434 n625 Dout_108 VDD GND NOR2_X1
xU12565 n8435 n628 Dout_111 VDD GND NOR2_X1
xU12566 n8435 n656 Dout_119 VDD GND NOR2_X1
xU12567 n8439 n188 Dout_0 VDD GND NOR2_X1
xU12568 n8436 n673 Dout_122 VDD GND NOR2_X1
xU12569 n8436 n301 Dout_16 VDD GND NOR2_X1
xU12570 n8439 n433 Dout_48 VDD GND NOR2_X1
xU12571 n8440 n459 Dout_56 VDD GND NOR2_X1
xU12572 n8440 n462 Dout_58 VDD GND NOR2_X1
xU12573 n8441 n483 Dout_64 VDD GND NOR2_X1
xU12574 n8443 n561 Dout_88 VDD GND NOR2_X1
xU12575 n8444 n570 Dout_93 VDD GND NOR2_X1
xU12576 n8434 n597 Dout_100 VDD GND NOR2_X1
xU12577 n8434 n617 Dout_104 VDD GND NOR2_X1
xU12578 n8434 n621 Dout_106 VDD GND NOR2_X1
xU12579 EN n137 VDD GND INV_X1
xU12580 n8437 n303 Dout_17 VDD GND NOR2_X1
xU12581 n8438 n388 Dout_33 VDD GND NOR2_X1
xU12582 n8440 n460 Dout_57 VDD GND NOR2_X1
xU12583 n8443 n539 Dout_81 VDD GND NOR2_X1
xU12584 n8436 n669 Dout_121 VDD GND NOR2_X1
xU12585 n8443 n563 Dout_89 VDD GND NOR2_X1
xU12586 n8437 n311 Dout_22 VDD GND NOR2_X1
xU12587 n8437 n312 Dout_23 VDD GND NOR2_X1
xU12588 n8440 n441 Dout_53 VDD GND NOR2_X1
xU12589 n8440 n443 Dout_55 VDD GND NOR2_X1
xU12590 n8442 n495 Dout_71 VDD GND NOR2_X1
xU12591 n8442 n519 Dout_78 VDD GND NOR2_X1
xU12592 n8444 n572 Dout_95 VDD GND NOR2_X1
xU12593 n8434 n600 Dout_103 VDD GND NOR2_X1
xU12594 n8434 n626 Dout_109 VDD GND NOR2_X1
xU12595 n8434 n248 Dout_10 VDD GND NOR2_X1
xU12596 n8436 n252 Dout_12 VDD GND NOR2_X1
xU12597 n8436 n254 Dout_14 VDD GND NOR2_X1
xU12598 n8437 n306 Dout_18 VDD GND NOR2_X1
xU12599 n8437 n361 Dout_24 VDD GND NOR2_X1
xU12600 n8438 n386 Dout_32 VDD GND NOR2_X1
xU12601 n8440 n436 Dout_50 VDD GND NOR2_X1
xU12602 n8444 n594 Dout_98 VDD GND NOR2_X1
xU12603 n8442 n513 Dout_73 VDD GND NOR2_X1
xU12604 n8442 n197 Dout_7 VDD GND NOR2_X1
xU12605 n8439 n418 Dout_47 VDD GND NOR2_X1
xU12606 n8443 n543 Dout_84 VDD GND NOR2_X1
xU12607 n8436 n678 Dout_125 VDD GND NOR2_X1
xU12608 n8438 n191 Dout_2 VDD GND NOR2_X1
xU12609 n8439 n415 Dout_44 VDD GND NOR2_X1
xU12610 n8442 n538 Dout_80 VDD GND NOR2_X1
xU12611 n8443 n541 Dout_82 VDD GND NOR2_X1
xU12612 n8435 n668 Dout_120 VDD GND NOR2_X1
xU12613 n8439 n411 Dout_41 VDD GND NOR2_X1
xU12614 n8437 n309 Dout_20 VDD GND NOR2_X1
xU12615 n8438 n368 Dout_30 VDD GND NOR2_X1
xU12616 n8438 n369 Dout_31 VDD GND NOR2_X1
xU12617 n8439 n395 Dout_39 VDD GND NOR2_X1
xU12618 n8440 n442 Dout_54 VDD GND NOR2_X1
xU12619 n8441 n466 Dout_61 VDD GND NOR2_X1
xU12620 n8441 n467 Dout_62 VDD GND NOR2_X1
xU12621 n8442 n494 Dout_70 VDD GND NOR2_X1
xU12622 n8444 n571 Dout_94 VDD GND NOR2_X1
xU12623 n8434 n598 Dout_101 VDD GND NOR2_X1
xU12624 n8435 n627 Dout_110 VDD GND NOR2_X1
xU12625 n8435 n647 Dout_113 VDD GND NOR2_X1
xU12626 n809 n7845 N3 VDD GND NOR2_X1
xU12627 Dvld_reg n8444 n7845 VDD GND OR2_X1
xU12628 n8436 n253 Dout_13 VDD GND NOR2_X1
xU12629 n8437 n310 Dout_21 VDD GND NOR2_X1
xU12630 n8437 n364 Dout_26 VDD GND NOR2_X1
xU12631 n8437 n365 Dout_27 VDD GND NOR2_X1
xU12632 n8438 n394 Dout_38 VDD GND NOR2_X1
xU12633 n8441 n489 Dout_66 VDD GND NOR2_X1
xU12634 n8442 n511 Dout_72 VDD GND NOR2_X1
xU12635 n8442 n515 Dout_74 VDD GND NOR2_X1
xU12636 n8442 n518 Dout_77 VDD GND NOR2_X1
xU12637 n8443 n565 Dout_90 VDD GND NOR2_X1
xU12638 n8443 n566 Dout_91 VDD GND NOR2_X1
xU12639 n8434 n599 Dout_102 VDD GND NOR2_X1
xU12640 n8435 n643 Dout_112 VDD GND NOR2_X1
xU12641 n8435 n650 Dout_114 VDD GND NOR2_X1
xU12642 n8435 n655 Dout_118 VDD GND NOR2_X1
xU12643 n8441 n195 Dout_5 VDD GND NOR2_X1
xU12644 n8441 n196 Dout_6 VDD GND NOR2_X1
xU12645 n8443 n544 Dout_85 VDD GND NOR2_X1
xU12646 n8443 n545 Dout_86 VDD GND NOR2_X1
xU12647 n8443 n546 Dout_87 VDD GND NOR2_X1
xU12648 n8436 n679 Dout_126 VDD GND NOR2_X1
xU12649 n8439 n417 Dout_46 VDD GND NOR2_X1
xU12650 n8439 n192 Dout_3 VDD GND NOR2_X1
xU12651 n8435 n249 Dout_11 VDD GND NOR2_X1
xU12652 n8437 n307 Dout_19 VDD GND NOR2_X1
xU12653 n8438 n389 Dout_34 VDD GND NOR2_X1
xU12654 n8438 n390 Dout_35 VDD GND NOR2_X1
xU12655 n8438 n393 Dout_37 VDD GND NOR2_X1
xU12656 n8439 n409 Dout_40 VDD GND NOR2_X1
xU12657 n8439 n412 Dout_42 VDD GND NOR2_X1
xU12658 n8439 n413 Dout_43 VDD GND NOR2_X1
xU12659 n8439 n416 Dout_45 VDD GND NOR2_X1
xU12660 n8440 n437 Dout_51 VDD GND NOR2_X1
xU12661 n8440 n463 Dout_59 VDD GND NOR2_X1
xU12662 n8441 n490 Dout_67 VDD GND NOR2_X1
xU12663 n8441 n493 Dout_69 VDD GND NOR2_X1
xU12664 n8442 n516 Dout_75 VDD GND NOR2_X1
xU12665 n8443 n542 Dout_83 VDD GND NOR2_X1
xU12666 n8434 n622 Dout_107 VDD GND NOR2_X1
xU12667 n8435 n651 Dout_115 VDD GND NOR2_X1
xU12668 n8435 n654 Dout_117 VDD GND NOR2_X1
xU12669 n8436 n674 Dout_123 VDD GND NOR2_X1
xU12670 n818 n7844 N4 VDD GND NOR2_X1
xU12671 n8444 Kvld_reg n7844 VDD GND OR2_X1
xU12672 n8444 n595 Dout_99 VDD GND NOR2_X1
xU12673 Kin_1 n127 VDD GND INV_X1
xU12674 Kin_104 n24 VDD GND INV_X1
xU12675 Kin_72 n56 VDD GND INV_X1
xU12676 Kin_112 n16 VDD GND INV_X1
xU12677 Kin_80 n48 VDD GND INV_X1
xU12678 Kin_120 n8 VDD GND INV_X1
xU12679 Kin_88 n40 VDD GND INV_X1
xU12680 Kin_96 n32 VDD GND INV_X1
xU12681 Kin_64 n64 VDD GND INV_X1
xU12682 Kin_32 n96 VDD GND INV_X1
xU12683 Kin_100 n28 VDD GND INV_X1
xU12684 Kin_68 n60 VDD GND INV_X1
xU12685 Kin_105 n23 VDD GND INV_X1
xU12686 Kin_73 n55 VDD GND INV_X1
xU12687 Kin_113 n15 VDD GND INV_X1
xU12688 Kin_81 n47 VDD GND INV_X1
xU12689 Kin_121 n7 VDD GND INV_X1
xU12690 Kin_89 n39 VDD GND INV_X1
xU12691 Kin_97 n31 VDD GND INV_X1
xU12692 Kin_65 n63 VDD GND INV_X1
xU12693 Kin_106 n22 VDD GND INV_X1
xU12694 Kin_74 n54 VDD GND INV_X1
xU12695 Kin_115 n13 VDD GND INV_X1
xU12696 Kin_83 n45 VDD GND INV_X1
xU12697 Kin_124 n4 VDD GND INV_X1
xU12698 Kin_92 n36 VDD GND INV_X1
xU12699 Kin_99 n29 VDD GND INV_X1
xU12700 Kin_67 n61 VDD GND INV_X1
xU12701 Kin_107 n21 VDD GND INV_X1
xU12702 Kin_75 n53 VDD GND INV_X1
xU12703 Kin_114 n14 VDD GND INV_X1
xU12704 Kin_82 n46 VDD GND INV_X1
xU12705 Kin_127 n1 VDD GND INV_X1
xU12706 Kin_95 n33 VDD GND INV_X1
xU12707 Kin_101 n27 VDD GND INV_X1
xU12708 Kin_69 n59 VDD GND INV_X1
xU12709 Kin_110 n18 VDD GND INV_X1
xU12710 Kin_78 n50 VDD GND INV_X1
xU12711 Kin_118 n10 VDD GND INV_X1
xU12712 Kin_86 n42 VDD GND INV_X1
xU12713 Kin_122 n6 VDD GND INV_X1
xU12714 Kin_90 n38 VDD GND INV_X1
xU12715 Kin_98 n30 VDD GND INV_X1
xU12716 Kin_66 n62 VDD GND INV_X1
xU12717 Kin_111 n17 VDD GND INV_X1
xU12718 Kin_79 n49 VDD GND INV_X1
xU12719 Kin_117 n11 VDD GND INV_X1
xU12720 Kin_85 n43 VDD GND INV_X1
xU12721 Kin_126 n2 VDD GND INV_X1
xU12722 Kin_94 n34 VDD GND INV_X1
xU12723 Kin_102 n26 VDD GND INV_X1
xU12724 Kin_70 n58 VDD GND INV_X1
xU12725 Kin_108 n20 VDD GND INV_X1
xU12726 Kin_76 n52 VDD GND INV_X1
xU12727 Kin_119 n9 VDD GND INV_X1
xU12728 Kin_87 n41 VDD GND INV_X1
xU12729 Kin_125 n3 VDD GND INV_X1
xU12730 Kin_93 n35 VDD GND INV_X1
xU12731 Kin_103 n25 VDD GND INV_X1
xU12732 Kin_71 n57 VDD GND INV_X1
xU12733 Kin_7 n121 VDD GND INV_X1
xU12734 Kin_39 n89 VDD GND INV_X1
xU12735 Kin_29 n99 VDD GND INV_X1
xU12736 Kin_61 n67 VDD GND INV_X1
xU12737 Kin_23 n105 VDD GND INV_X1
xU12738 Kin_55 n73 VDD GND INV_X1
xU12739 Kin_116 n12 VDD GND INV_X1
xU12740 Kin_84 n44 VDD GND INV_X1
xU12741 Kin_20 n108 VDD GND INV_X1
xU12742 Kin_52 n76 VDD GND INV_X1
xU12743 Kin_12 n116 VDD GND INV_X1
xU12744 Kin_44 n84 VDD GND INV_X1
xU12745 Kin_6 n122 VDD GND INV_X1
xU12746 Kin_38 n90 VDD GND INV_X1
xU12747 Kin_30 n98 VDD GND INV_X1
xU12748 Kin_62 n66 VDD GND INV_X1
xU12749 Kin_21 n107 VDD GND INV_X1
xU12750 Kin_53 n75 VDD GND INV_X1
xU12751 Kin_15 n113 VDD GND INV_X1
xU12752 Kin_47 n81 VDD GND INV_X1
xU12753 Kin_2 n126 VDD GND INV_X1
xU12754 Kin_34 n94 VDD GND INV_X1
xU12755 Kin_26 n102 VDD GND INV_X1
xU12756 Kin_58 n70 VDD GND INV_X1
xU12757 Kin_22 n106 VDD GND INV_X1
xU12758 Kin_54 n74 VDD GND INV_X1
xU12759 Kin_14 n114 VDD GND INV_X1
xU12760 Kin_46 n82 VDD GND INV_X1
xU12761 Kin_5 n123 VDD GND INV_X1
xU12762 Kin_37 n91 VDD GND INV_X1
xU12763 Kin_31 n97 VDD GND INV_X1
xU12764 Kin_63 n65 VDD GND INV_X1
xU12765 Kin_18 n110 VDD GND INV_X1
xU12766 Kin_50 n78 VDD GND INV_X1
xU12767 Kin_11 n117 VDD GND INV_X1
xU12768 Kin_43 n85 VDD GND INV_X1
xU12769 Kin_109 n19 VDD GND INV_X1
xU12770 Kin_77 n51 VDD GND INV_X1
xU12771 Kin_13 n115 VDD GND INV_X1
xU12772 Kin_45 n83 VDD GND INV_X1
xU12773 Kin_3 n125 VDD GND INV_X1
xU12774 Kin_35 n93 VDD GND INV_X1
xU12775 Kin_28 n100 VDD GND INV_X1
xU12776 Kin_60 n68 VDD GND INV_X1
xU12777 Kin_123 n5 VDD GND INV_X1
xU12778 Kin_91 n37 VDD GND INV_X1
xU12779 Kin_27 n101 VDD GND INV_X1
xU12780 Kin_59 n69 VDD GND INV_X1
xU12781 Kin_19 n109 VDD GND INV_X1
xU12782 Kin_51 n77 VDD GND INV_X1
xU12783 Kin_10 n118 VDD GND INV_X1
xU12784 Kin_42 n86 VDD GND INV_X1
xU12785 Kin_33 n95 VDD GND INV_X1
xU12786 Kin_25 n103 VDD GND INV_X1
xU12787 Kin_57 n71 VDD GND INV_X1
xU12788 Kin_17 n111 VDD GND INV_X1
xU12789 Kin_49 n79 VDD GND INV_X1
xU12790 Kin_9 n119 VDD GND INV_X1
xU12791 Kin_41 n87 VDD GND INV_X1
xU12792 Kin_4 n124 VDD GND INV_X1
xU12793 Kin_36 n92 VDD GND INV_X1
xU12794 Kin_24 n104 VDD GND INV_X1
xU12795 Kin_56 n72 VDD GND INV_X1
xU12796 Kin_16 n112 VDD GND INV_X1
xU12797 Kin_48 n80 VDD GND INV_X1
xU12798 Kin_8 n120 VDD GND INV_X1
xU12799 Kin_40 n88 VDD GND INV_X1
xU12800 Kin_0 n128 VDD GND INV_X1
xU12801 n8271 n8281 VDD GND INV_X1
xU12802 n8282 n8291 VDD GND BUF_X1
xU12803 n8282 n8292 VDD GND BUF_X1
xU12804 n8282 n8293 VDD GND BUF_X1
xU12805 n8282 n8294 VDD GND BUF_X1
xU12806 n8282 n8295 VDD GND BUF_X1
xU12807 n8283 n8296 VDD GND BUF_X1
xU12808 n8283 n8297 VDD GND BUF_X1
xU12809 n8283 n8298 VDD GND BUF_X1
xU12810 n8283 n8299 VDD GND BUF_X1
xU12811 n8283 n8300 VDD GND BUF_X1
xU12812 n8284 n8301 VDD GND BUF_X1
xU12813 n8284 n8302 VDD GND BUF_X1
xU12814 n8284 n8303 VDD GND BUF_X1
xU12815 n8284 n8304 VDD GND BUF_X1
xU12816 n8284 n8305 VDD GND BUF_X1
xU12817 n8285 n8306 VDD GND BUF_X1
xU12818 n8285 n8307 VDD GND BUF_X1
xU12819 n8285 n8308 VDD GND BUF_X1
xU12820 n8285 n8309 VDD GND BUF_X1
xU12821 n8340 n8326 VDD GND INV_X1
xU12822 n8340 n8327 VDD GND INV_X1
xU12823 n8340 n8328 VDD GND INV_X1
xU12824 n1009 n8341 VDD GND BUF_X1
xU12825 n1009 n8342 VDD GND BUF_X1
xU12826 n1009 n8343 VDD GND BUF_X1
xU12827 n1009 n8344 VDD GND BUF_X1
xU12828 n1009 n8345 VDD GND BUF_X1
xU12829 n1009 n8351 VDD GND BUF_X1
xU12830 n1007 n8352 VDD GND BUF_X1
xU12831 n1007 n8353 VDD GND BUF_X1
xU12832 n1007 n8354 VDD GND BUF_X1
xU12833 n1007 n8355 VDD GND BUF_X1
xU12834 n1007 n8356 VDD GND BUF_X1
xU12835 n8356 n8370 VDD GND BUF_X1
xU12836 n991 n8371 VDD GND BUF_X1
xU12837 n991 n8372 VDD GND BUF_X1
xU12838 n991 n8373 VDD GND BUF_X1
xU12839 n991 n8374 VDD GND BUF_X1
xU12840 n991 n8375 VDD GND BUF_X1
xU12841 n991 n8376 VDD GND BUF_X1
xU12842 n991 n8377 VDD GND BUF_X1
xU12843 n8377 n8398 VDD GND BUF_X1
xU12844 n8399 n8402 VDD GND BUF_X1
xU12845 n8399 n8403 VDD GND BUF_X1
xU12846 n8399 n8404 VDD GND BUF_X1
xU12847 n8399 n8405 VDD GND BUF_X1
xU12848 n8399 n8406 VDD GND BUF_X1
xU12849 n8399 n8407 VDD GND BUF_X1
xU12850 n8400 n8413 VDD GND BUF_X1
xU12851 n8400 n8414 VDD GND BUF_X1
xU12852 n8400 n8415 VDD GND BUF_X1
xU12853 n8400 n8416 VDD GND BUF_X1
xU12854 n8400 n8417 VDD GND BUF_X1
xU12855 n8400 n8418 VDD GND BUF_X1
xU12856 n8401 n8424 VDD GND BUF_X1
xU12857 n8401 n8425 VDD GND BUF_X1
xU12858 n8401 n8426 VDD GND BUF_X1
xU12859 n8401 n8427 VDD GND BUF_X1
xU12860 n8401 n8433 VDD GND BUF_X1



.PRINT TRAN V(N3) V(VDD)

.END
