.Option ingold=2 accurate
.OPTION MEASDGT=8
.OPTION NUMDGT=10
+ RUNLVL=5 ACCURATE
.op
.PARAM LMIN='50E-9'
.PARAM VDD_VALUE= 1.2
.PARAM VDD_HALF= 0.6
.OPTION BRIEF=1

.OPTION POST=2
.OPTION MEASFORM=3
.OPTION PROBE=1

VSUPPLY VDD 0 VDD_VALUE
VSUPPLYGND GND 0 0

Vinput CLK GND PULSE(0 1.2 0.0001n 0.0001n 0.0001n .2465n .495n)
*Vclk CLK GND PULSE(0 1.2 0.0001n 0.0001n 0.0001n 0.33n .66n)
*PULSE (v1 v2 <td <tr <tf <pw <per>>>>>)

.TRAN .2475N 25N START=0N

.include './trans_model_nk'
.temp 0

******** NAND MODEL ***********
* The subcircuit for NAND
.SUBCKT NAND2_X1
+ A1 A2
+ ZN
+ VDDx GNDx
M_i_1 net_0 A1 GNDx GNDx NMOS_VTL W=0.415000U L='LMIN'
M_i_0 ZN A2 net_0 GNDx NMOS_VTL W=0.415000U L='LMIN'
M_i_11 ZN A2 VDDx VDDx PMOS_VTL W=0.630000U L='LMIN'
M_i_10 VDDx A1 ZN VDDx PMOS_VTL W=0.630000U L='LMIN'
.ENDS

******** INV MODEL ***********
* The subcircuit for INV
.SUBCKT INV_X1
+ A1
+ ZN
+ VDDx GNDx
M_i_0 ZN A1 GNDx GNDx NMOS_VTL W=0.415000U L='LMIN'
M_i_10 ZN A1 VDDx VDDx PMOS_VTL W=0.630000U L='LMIN'
.ENDS

******** DFFR_X1 MODEL ***********
* The subcircuit for DFFR_X1
.SUBCKT DFFR_X1
+ D CK RN
+ Q QN
+ VDDx GNDx

*.PININFO D:I RN:I CK:I Q:O QN:O VDDx:P GNDx:G 
M_i_0 GNDx CK net_000 GNDx NMOS_VTL W=0.210000U L='LMIN'
M_i_7 net_001 net_000 GNDx GNDx NMOS_VTL W=0.210000U L='LMIN'
M_i_13 net_002 D GNDx GNDx NMOS_VTL W=0.275000U L='LMIN'
M_i_18 net_003 net_000 net_002 GNDx NMOS_VTL W=0.275000U L='LMIN'
M_i_24 net_004 net_001 net_003 GNDx NMOS_VTL W=0.090000U L='LMIN'
M_i_28 net_005 net_006 net_004 GNDx NMOS_VTL W=0.090000U L='LMIN'
M_i_32 GNDx RN net_005 GNDx NMOS_VTL W=0.090000U L='LMIN'
M_i_38 GNDx net_003 net_006 GNDx NMOS_VTL W=0.210000U L='LMIN'
M_i_45 net_007 net_003 GNDx GNDx NMOS_VTL W=0.210000U L='LMIN'
M_i_49 net_008 net_001 net_007 GNDx NMOS_VTL W=0.210000U L='LMIN'
M_i_55 net_009 net_000 net_008 GNDx NMOS_VTL W=0.090000U L='LMIN'
M_i_59 GNDx net_011 net_009 GNDx NMOS_VTL W=0.090000U L='LMIN'
M_i_65 net_010 RN GNDx GNDx NMOS_VTL W=0.210000U L='LMIN'
M_i_70 net_011 net_008 net_010 GNDx NMOS_VTL W=0.210000U L='LMIN'
M_i_76 GNDx net_008 QN GNDx NMOS_VTL W=0.415000U L='LMIN'
M_i_83 Q net_011 GNDx GNDx NMOS_VTL W=0.415000U L='LMIN'
M_i_89 VDDx CK net_000 VDDx PMOS_VTL W=0.315000U L='LMIN'
M_i_96 net_001 net_000 VDDx VDDx PMOS_VTL W=0.315000U L='LMIN'
M_i_103 net_012 D VDDx VDDx PMOS_VTL W=0.420000U L='LMIN'
M_i_108 net_003 net_001 net_012 VDDx PMOS_VTL W=0.420000U L='LMIN'
M_i_114 net_013 net_000 net_003 VDDx PMOS_VTL W=0.090000U L='LMIN'
M_i_119 VDDx net_006 net_013 VDDx PMOS_VTL W=0.090000U L='LMIN'
M_i_125 net_013 RN VDDx VDDx PMOS_VTL W=0.090000U L='LMIN'
M_i_136 VDDx net_003 net_006 VDDx PMOS_VTL W=0.315000U L='LMIN'
M_i_143 net_015 net_003 VDDx VDDx PMOS_VTL W=0.315000U L='LMIN'
M_i_147 net_008 net_000 net_015 VDDx PMOS_VTL W=0.315000U L='LMIN'
M_i_153 net_016 net_001 net_008 VDDx PMOS_VTL W=0.090000U L='LMIN'
M_i_159 VDDx net_011 net_016 VDDx PMOS_VTL W=0.090000U L='LMIN'
M_i_165 net_011 RN VDDx VDDx PMOS_VTL W=0.315000U L='LMIN'
M_i_172 VDDx net_008 net_011 VDDx PMOS_VTL W=0.315000U L='LMIN'
M_i_180 VDDx net_008 QN VDDx PMOS_VTL W=0.630000U L='LMIN'
M_i_187 Q net_011 VDDx VDDx PMOS_VTL W=0.630000U L='LMIN'
.ENDS 

**Ringoscillator
XNand1 A1 A2 ZN VDD GND NAND2_X1

Xinv2 A1 ZN VDD GND INV_X1
Xinv3 A1 ZN VDD GND INV_X1
Xinv4 A1 ZN VDD GND INV_X1
Xinv5 A1 ZN VDD GND INV_X1
Xinv6 A1 ZN VDD GND INV_X1
Xinv7 A1 ZN VDD GND INV_X1
Xinv8 A1 ZN VDD GND INV_X1
Xinv9 A1 ZN VDD GND INV_X1
Xinv10 A1 ZN VDD GND INV_X1
Xinv11 A1 ZN VDD GND INV_X1
Xinv12 A1 ZN VDD GND INV_X1
Xinv13 A1 ZN VDD GND INV_X1
Xinv14 A1 ZN VDD GND INV_X1
Xinv15 A1 ZN VDD GND INV_X1
Xinv16 A1 ZN VDD GND INV_X1
Xinv17 A1 ZN VDD GND INV_X1
Xinv18 A1 ZN VDD GND INV_X1
Xinv19 A1 ZN VDD GND INV_X1
Xinv20 A1 ZN VDD GND INV_X1
Xinv21 A1 ZN VDD GND INV_X1

**Counter

XDFF0 CK RN Q QN VDD GND DFFR_X1
XDFF1 CK RN Q QN VDD GND DFFR_X1
XDFF2 CK RN Q QN VDD GND DFFR_X1
XDFF3 CK RN Q QN VDD GND DFFR_X1
XDFF4 CK RN Q QN VDD GND DFFR_X1
XDFF5 CK RN Q QN VDD GND DFFR_X1
XDFF6 CK RN Q QN VDD GND DFFR_X1
XDFF7 CK RN Q QN VDD GND DFFR_X1
XDFF8 CK RN Q QN VDD GND DFFR_X1
XDFF9 CK RN Q QN VDD GND DFFR_X1
    


* The monitoring
.PRINT TRAN 


.END