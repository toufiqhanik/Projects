`timescale 1ns / 1ps


module softbox(din, dout);

input [7:0] din;
output [7:0] dout;

reg [7:0] sv;


always @(din)
    case (din)

       8'h00: sv=8'h63;
	   8'h01: sv=8'h7c;
	   8'h02: sv=8'h77;
	   8'h03: sv=8'h7b;
	   8'h04: sv=8'hf2;
	   8'h05: sv=8'h6b;
	   8'h06: sv=8'h6f;
	   8'h07: sv=8'hc5;
	   8'h08: sv=8'h30;
	   8'h09: sv=8'h01;
	   8'h0a: sv=8'h67;
	   8'h0b: sv=8'h2b;
	   8'h0c: sv=8'hfe;
	   8'h0d: sv=8'hd7;
	   8'h0e: sv=8'hab;
	   8'h0f: sv=8'h76;
	   8'h10: sv=8'hca;
	   8'h11: sv=8'h82;
	   8'h12: sv=8'hc9;
	   8'h13: sv=8'h7d;
	   8'h14: sv=8'hfa;
	   8'h15: sv=8'h59;
	   8'h16: sv=8'h47;
	   8'h17: sv=8'hf0;
	   8'h18: sv=8'had;
	   8'h19: sv=8'hd4;
	   8'h1a: sv=8'ha2;
	   8'h1b: sv=8'haf;
	   8'h1c: sv=8'h9c;
	   8'h1d: sv=8'ha4;
	   8'h1e: sv=8'h72;
	   8'h1f: sv=8'hc0;
	   8'h20: sv=8'hb7;
	   8'h21: sv=8'hfd;
	   8'h22: sv=8'h93;
	   8'h23: sv=8'h26;
	   8'h24: sv=8'h36;
	   8'h25: sv=8'h3f;
	   8'h26: sv=8'hf7;
	   8'h27: sv=8'hcc;
	   8'h28: sv=8'h34;
	   8'h29: sv=8'ha5;
	   8'h2a: sv=8'he5;
	   8'h2b: sv=8'hf1;
	   8'h2c: sv=8'h71;
	   8'h2d: sv=8'hd8;
	   8'h2e: sv=8'h31;
	   8'h2f: sv=8'h15;
	   8'h30: sv=8'h04;
	   8'h31: sv=8'hc7;
	   8'h32: sv=8'h23;
	   8'h33: sv=8'hc3;
	   8'h34: sv=8'h18;
	   8'h35: sv=8'h96;
	   8'h36: sv=8'h05;
	   8'h37: sv=8'h9a;
	   8'h38: sv=8'h07;
	   8'h39: sv=8'h12;
	   8'h3a: sv=8'h80;
	   8'h3b: sv=8'he2;
	   8'h3c: sv=8'heb;
	   8'h3d: sv=8'h27;
	   8'h3e: sv=8'hb2;
	   8'h3f: sv=8'h75;
	   8'h40: sv=8'h09;
	   8'h41: sv=8'h83;
	   8'h42: sv=8'h2c;
	   8'h43: sv=8'h1a;
	   8'h44: sv=8'h1b;
	   8'h45: sv=8'h6e;
	   8'h46: sv=8'h5a;
	   8'h47: sv=8'ha0;
	   8'h48: sv=8'h52;
	   8'h49: sv=8'h3b;
	   8'h4a: sv=8'hd6;
	   8'h4b: sv=8'hb3;
	   8'h4c: sv=8'h29;
	   8'h4d: sv=8'he3;
	   8'h4e: sv=8'h2f;
	   8'h4f: sv=8'h84;
	   8'h50: sv=8'h53;
	   8'h51: sv=8'hd1;
	   8'h52: sv=8'h00;
	   8'h53: sv=8'hed;
	   8'h54: sv=8'h20;
	   8'h55: sv=8'hfc;
	   8'h56: sv=8'hb1;
	   8'h57: sv=8'h5b;
	   8'h58: sv=8'h6a;
	   8'h59: sv=8'hcb;
	   8'h5a: sv=8'hbe;
	   8'h5b: sv=8'h39;
	   8'h5c: sv=8'h4a;
	   8'h5d: sv=8'h4c;
	   8'h5e: sv=8'h58;
	   8'h5f: sv=8'hcf;
	   8'h60: sv=8'hd0;
	   8'h61: sv=8'hef;
	   8'h62: sv=8'haa;
	   8'h63: sv=8'hfb;
	   8'h64: sv=8'h43;
	   8'h65: sv=8'h4d;
	   8'h66: sv=8'h33;
	   8'h67: sv=8'h85;
	   8'h68: sv=8'h45;
	   8'h69: sv=8'hf9;
	   8'h6a: sv=8'h02;
	   8'h6b: sv=8'h7f;
	   8'h6c: sv=8'h50;
	   8'h6d: sv=8'h3c;
	   8'h6e: sv=8'h9f;
	   8'h6f: sv=8'ha8;
	   8'h70: sv=8'h51;
	   8'h71: sv=8'ha3;
	   8'h72: sv=8'h40;
	   8'h73: sv=8'h8f;
	   8'h74: sv=8'h92;
	   8'h75: sv=8'h9d;
	   8'h76: sv=8'h38;
	   8'h77: sv=8'hf5;
	   8'h78: sv=8'hbc;
	   8'h79: sv=8'hb6;
	   8'h7a: sv=8'hda;
	   8'h7b: sv=8'h21;
	   8'h7c: sv=8'h10;
	   8'h7d: sv=8'hff;
	   8'h7e: sv=8'hf3;
	   8'h7f: sv=8'hd2;
	   8'h80: sv=8'hcd;
	   8'h81: sv=8'h0c;
	   8'h82: sv=8'h13;
	   8'h83: sv=8'hec;
	   8'h84: sv=8'h5f;
	   8'h85: sv=8'h97;
	   8'h86: sv=8'h44;
	   8'h87: sv=8'h17;
	   8'h88: sv=8'hc4;
	   8'h89: sv=8'ha7;
	   8'h8a: sv=8'h7e;
	   8'h8b: sv=8'h3d;
	   8'h8c: sv=8'h64;
	   8'h8d: sv=8'h5d;
	   8'h8e: sv=8'h19;
	   8'h8f: sv=8'h73;
	   8'h90: sv=8'h60;
	   8'h91: sv=8'h81;
	   8'h92: sv=8'h4f;
	   8'h93: sv=8'hdc;
	   8'h94: sv=8'h22;
	   8'h95: sv=8'h2a;
	   8'h96: sv=8'h90;
	   8'h97: sv=8'h88;
	   8'h98: sv=8'h46;
	   8'h99: sv=8'hee;
	   8'h9a: sv=8'hb8;
	   8'h9b: sv=8'h14;
	   8'h9c: sv=8'hde;
	   8'h9d: sv=8'h5e;
	   8'h9e: sv=8'h0b;
	   8'h9f: sv=8'hdb;
	   8'ha0: sv=8'he0;
	   8'ha1: sv=8'h32;
	   8'ha2: sv=8'h3a;
	   8'ha3: sv=8'h0a;
	   8'ha4: sv=8'h49;
	   8'ha5: sv=8'h06;
	   8'ha6: sv=8'h24;
	   8'ha7: sv=8'h5c;
	   8'ha8: sv=8'hc2;
	   8'ha9: sv=8'hd3;
	   8'haa: sv=8'hac;
	   8'hab: sv=8'h62;
	   8'hac: sv=8'h91;
	   8'had: sv=8'h95;
	   8'hae: sv=8'he4;
	   8'haf: sv=8'h79;
	   8'hb0: sv=8'he7;
	   8'hb1: sv=8'hc8;
	   8'hb2: sv=8'h37;
	   8'hb3: sv=8'h6d;
	   8'hb4: sv=8'h8d;
	   8'hb5: sv=8'hd5;
	   8'hb6: sv=8'h4e;
	   8'hb7: sv=8'ha9;
	   8'hb8: sv=8'h6c;
	   8'hb9: sv=8'h56;
	   8'hba: sv=8'hf4;
	   8'hbb: sv=8'hea;
	   8'hbc: sv=8'h65;
	   8'hbd: sv=8'h7a;
	   8'hbe: sv=8'hae;
	   8'hbf: sv=8'h08;
	   8'hc0: sv=8'hba;
	   8'hc1: sv=8'h78;
	   8'hc2: sv=8'h25;
	   8'hc3: sv=8'h2e;
	   8'hc4: sv=8'h1c;
	   8'hc5: sv=8'ha6;
	   8'hc6: sv=8'hb4;
	   8'hc7: sv=8'hc6;
	   8'hc8: sv=8'he8;
	   8'hc9: sv=8'hdd;
	   8'hca: sv=8'h74;
	   8'hcb: sv=8'h1f;
	   8'hcc: sv=8'h4b;
	   8'hcd: sv=8'hbd;
	   8'hce: sv=8'h8b;
	   8'hcf: sv=8'h8a;
	   8'hd0: sv=8'h70;
	   8'hd1: sv=8'h3e;
	   8'hd2: sv=8'hb5;
	   8'hd3: sv=8'h66;
	   8'hd4: sv=8'h48;
	   8'hd5: sv=8'h03;
	   8'hd6: sv=8'hf6;
	   8'hd7: sv=8'h0e;
	   8'hd8: sv=8'h61;
	   8'hd9: sv=8'h35;
	   8'hda: sv=8'h57;
	   8'hdb: sv=8'hb9;
	   8'hdc: sv=8'h86;
	   8'hdd: sv=8'hc1;
	   8'hde: sv=8'h1d;
	   8'hdf: sv=8'h9e;
	   8'he0: sv=8'he1;
	   8'he1: sv=8'hf8;
	   8'he2: sv=8'h98;
	   8'he3: sv=8'h11;
	   8'he4: sv=8'h69;
	   8'he5: sv=8'hd9;
	   8'he6: sv=8'h8e;
	   8'he7: sv=8'h94;
	   8'he8: sv=8'h9b;
	   8'he9: sv=8'h1e;
	   8'hea: sv=8'h87;
	   8'heb: sv=8'he9;
	   8'hec: sv=8'hce;
	   8'hed: sv=8'h55;
	   8'hee: sv=8'h28;
	   8'hef: sv=8'hdf;
	   8'hf0: sv=8'h8c;
	   8'hf1: sv=8'ha1;
	   8'hf2: sv=8'h89;
	   8'hf3: sv=8'h0d;
	   8'hf4: sv=8'hbf;
	   8'hf5: sv=8'he6;
	   8'hf6: sv=8'h42;
	   8'hf7: sv=8'h68;
	   8'hf8: sv=8'h41;
	   8'hf9: sv=8'h99;
	   8'hfa: sv=8'h2d;
	   8'hfb: sv=8'h0f;
	   8'hfc: sv=8'hb0;
	   8'hfd: sv=8'h54;
	   8'hfe: sv=8'hbb;
	   8'hff: sv=8'h16;
	endcase

	assign dout = sv;

endmodule

